`timescale 1ns / 1ps

module ann_weights_and_biases();

parameter WEIGHT_0_0 = 16'd-1836;
parameter WEIGHT_0_1 = 16'd-720;
parameter WEIGHT_0_2 = 16'd-977;
parameter WEIGHT_0_3 = 16'd-2697;
parameter WEIGHT_0_4 = 16'd2430;
parameter WEIGHT_0_5 = 16'd1817;
parameter WEIGHT_0_6 = 16'd1425;
parameter WEIGHT_0_7 = 16'd1812;
parameter WEIGHT_0_8 = 16'd-1636;
parameter WEIGHT_0_9 = 16'd833;
parameter WEIGHT_0_10 = 16'd-1022;
parameter WEIGHT_0_11 = 16'd164;
parameter WEIGHT_0_12 = 16'd-1184;
parameter WEIGHT_0_13 = 16'd1665;
parameter WEIGHT_0_14 = 16'd-590;
parameter WEIGHT_0_15 = 16'd1614;
parameter WEIGHT_0_16 = 16'd720;
parameter WEIGHT_0_17 = 16'd-1761;
parameter WEIGHT_0_18 = 16'd2372;
parameter WEIGHT_0_19 = 16'd-2446;
parameter WEIGHT_0_20 = 16'd2223;
parameter WEIGHT_0_21 = 16'd-2314;
parameter WEIGHT_0_22 = 16'd-1300;
parameter WEIGHT_0_23 = 16'd-1179;
parameter WEIGHT_0_24 = 16'd-161;
parameter WEIGHT_0_25 = 16'd2447;
parameter WEIGHT_0_26 = 16'd-2403;
parameter WEIGHT_0_27 = 16'd2258;
parameter WEIGHT_0_28 = 16'd2629;
parameter WEIGHT_0_29 = 16'd1415;
parameter WEIGHT_0_30 = 16'd85;
parameter WEIGHT_0_31 = 16'd-680;
parameter WEIGHT_0_32 = 16'd-1705;
parameter WEIGHT_0_33 = 16'd145;
parameter WEIGHT_0_34 = 16'd310;
parameter WEIGHT_0_35 = 16'd-2751;
parameter WEIGHT_0_36 = 16'd-2376;
parameter WEIGHT_0_37 = 16'd-863;
parameter WEIGHT_0_38 = 16'd2469;
parameter WEIGHT_0_39 = 16'd1513;
parameter WEIGHT_0_40 = 16'd-702;
parameter WEIGHT_0_41 = 16'd704;
parameter WEIGHT_0_42 = 16'd458;
parameter WEIGHT_0_43 = 16'd-707;
parameter WEIGHT_0_44 = 16'd-2805;
parameter WEIGHT_0_45 = 16'd-1317;
parameter WEIGHT_0_46 = 16'd-1795;
parameter WEIGHT_0_47 = 16'd-1651;
parameter WEIGHT_0_48 = 16'd641;
parameter WEIGHT_0_49 = 16'd-767;
parameter WEIGHT_0_50 = 16'd-719;
parameter WEIGHT_0_51 = 16'd1880;
parameter WEIGHT_0_52 = 16'd2668;
parameter WEIGHT_0_53 = 16'd-1678;
parameter WEIGHT_0_54 = 16'd2240;
parameter WEIGHT_0_55 = 16'd-2530;
parameter WEIGHT_0_56 = 16'd1017;
parameter WEIGHT_0_57 = 16'd612;
parameter WEIGHT_0_58 = 16'd1967;
parameter WEIGHT_0_59 = 16'd-1244;
parameter WEIGHT_0_60 = 16'd-2742;
parameter WEIGHT_0_61 = 16'd-1157;
parameter WEIGHT_0_62 = 16'd-2383;
parameter WEIGHT_0_63 = 16'd-2670;
parameter WEIGHT_0_64 = 16'd1583;
parameter WEIGHT_0_65 = 16'd-2479;
parameter WEIGHT_0_66 = 16'd180;
parameter WEIGHT_0_67 = 16'd2656;
parameter WEIGHT_0_68 = 16'd2079;
parameter WEIGHT_0_69 = 16'd2826;
parameter WEIGHT_0_70 = 16'd-2106;
parameter WEIGHT_0_71 = 16'd-881;
parameter WEIGHT_0_72 = 16'd-173;
parameter WEIGHT_0_73 = 16'd158;
parameter WEIGHT_0_74 = 16'd-288;
parameter WEIGHT_0_75 = 16'd-627;
parameter WEIGHT_0_76 = 16'd-985;
parameter WEIGHT_0_77 = 16'd-1543;
parameter WEIGHT_0_78 = 16'd-1641;
parameter WEIGHT_0_79 = 16'd-2283;
parameter WEIGHT_0_80 = 16'd-1895;
parameter WEIGHT_0_81 = 16'd1757;
parameter WEIGHT_0_82 = 16'd350;
parameter WEIGHT_0_83 = 16'd24;
parameter WEIGHT_0_84 = 16'd14;
parameter WEIGHT_0_85 = 16'd397;
parameter WEIGHT_0_86 = 16'd-1989;
parameter WEIGHT_0_87 = 16'd-1952;
parameter WEIGHT_0_88 = 16'd-228;
parameter WEIGHT_0_89 = 16'd-49;
parameter WEIGHT_0_90 = 16'd1836;
parameter WEIGHT_0_91 = 16'd853;
parameter WEIGHT_0_92 = 16'd-1136;
parameter WEIGHT_0_93 = 16'd747;
parameter WEIGHT_0_94 = 16'd-1314;
parameter WEIGHT_0_95 = 16'd-1347;
parameter WEIGHT_0_96 = 16'd-2015;
parameter WEIGHT_0_97 = 16'd2724;
parameter WEIGHT_0_98 = 16'd1334;
parameter WEIGHT_0_99 = 16'd1197;
parameter WEIGHT_0_100 = 16'd-1449;
parameter WEIGHT_0_101 = 16'd-2673;
parameter WEIGHT_0_102 = 16'd1157;
parameter WEIGHT_0_103 = 16'd2531;
parameter WEIGHT_0_104 = 16'd-168;
parameter WEIGHT_0_105 = 16'd100;
parameter WEIGHT_0_106 = 16'd2168;
parameter WEIGHT_0_107 = 16'd-2204;
parameter WEIGHT_0_108 = 16'd2292;
parameter WEIGHT_0_109 = 16'd1555;
parameter WEIGHT_0_110 = 16'd-961;
parameter WEIGHT_0_111 = 16'd-1483;
parameter WEIGHT_0_112 = 16'd2550;
parameter WEIGHT_0_113 = 16'd2258;
parameter WEIGHT_0_114 = 16'd-2132;
parameter WEIGHT_0_115 = 16'd1923;
parameter WEIGHT_0_116 = 16'd2049;
parameter WEIGHT_0_117 = 16'd2132;
parameter WEIGHT_0_118 = 16'd-28;
parameter WEIGHT_0_119 = 16'd138;
parameter WEIGHT_0_120 = 16'd-2588;
parameter WEIGHT_0_121 = 16'd-33;
parameter WEIGHT_0_122 = 16'd-2350;
parameter WEIGHT_0_123 = 16'd-2339;
parameter WEIGHT_0_124 = 16'd-3578;
parameter WEIGHT_0_125 = 16'd-678;
parameter WEIGHT_0_126 = 16'd883;
parameter WEIGHT_0_127 = 16'd-970;
parameter WEIGHT_0_128 = 16'd-2418;
parameter WEIGHT_0_129 = 16'd-3801;
parameter WEIGHT_0_130 = 16'd-1548;
parameter WEIGHT_0_131 = 16'd-2588;
parameter WEIGHT_0_132 = 16'd1053;
parameter WEIGHT_0_133 = 16'd-5012;
parameter WEIGHT_0_134 = 16'd-568;
parameter WEIGHT_0_135 = 16'd-3308;
parameter WEIGHT_0_136 = 16'd4781;
parameter WEIGHT_0_137 = 16'd69;
parameter WEIGHT_0_138 = 16'd-4880;
parameter WEIGHT_0_139 = 16'd-2167;
parameter WEIGHT_0_140 = 16'd-3039;
parameter WEIGHT_0_141 = 16'd-2506;
parameter WEIGHT_0_142 = 16'd3585;
parameter WEIGHT_0_143 = 16'd-647;
parameter WEIGHT_0_144 = 16'd-3209;
parameter WEIGHT_0_145 = 16'd409;
parameter WEIGHT_0_146 = 16'd-2512;
parameter WEIGHT_0_147 = 16'd-1752;
parameter WEIGHT_0_148 = 16'd1252;
parameter WEIGHT_0_149 = 16'd-3695;
parameter WEIGHT_0_150 = 16'd-655;
parameter WEIGHT_0_151 = 16'd-1990;
parameter WEIGHT_0_152 = 16'd942;
parameter WEIGHT_0_153 = 16'd-2595;
parameter WEIGHT_0_154 = 16'd-3623;
parameter WEIGHT_0_155 = 16'd1213;
parameter WEIGHT_0_156 = 16'd699;
parameter WEIGHT_0_157 = 16'd-1394;
parameter WEIGHT_0_158 = 16'd-2593;
parameter WEIGHT_0_159 = 16'd-1423;
parameter WEIGHT_0_160 = 16'd2622;
parameter WEIGHT_0_161 = 16'd-1094;
parameter WEIGHT_0_162 = 16'd-74;
parameter WEIGHT_0_163 = 16'd-171;
parameter WEIGHT_0_164 = 16'd-2311;
parameter WEIGHT_0_165 = 16'd-2478;
parameter WEIGHT_0_166 = 16'd-1896;
parameter WEIGHT_0_167 = 16'd-1610;
parameter WEIGHT_0_168 = 16'd-1411;
parameter WEIGHT_0_169 = 16'd-318;
parameter WEIGHT_0_170 = 16'd-1210;
parameter WEIGHT_0_171 = 16'd1450;
parameter WEIGHT_0_172 = 16'd-519;
parameter WEIGHT_0_173 = 16'd1886;
parameter WEIGHT_0_174 = 16'd2492;
parameter WEIGHT_0_175 = 16'd481;
parameter WEIGHT_0_176 = 16'd134;
parameter WEIGHT_0_177 = 16'd109;
parameter WEIGHT_0_178 = 16'd-724;
parameter WEIGHT_0_179 = 16'd-2690;
parameter WEIGHT_0_180 = 16'd2365;
parameter WEIGHT_0_181 = 16'd-2609;
parameter WEIGHT_0_182 = 16'd-1421;
parameter WEIGHT_0_183 = 16'd2456;
parameter WEIGHT_0_184 = 16'd-980;
parameter WEIGHT_0_185 = 16'd-509;
parameter WEIGHT_0_186 = 16'd1844;
parameter WEIGHT_0_187 = 16'd308;
parameter WEIGHT_0_188 = 16'd-1455;
parameter WEIGHT_0_189 = 16'd495;
parameter WEIGHT_0_190 = 16'd2239;
parameter WEIGHT_0_191 = 16'd2273;
parameter WEIGHT_0_192 = 16'd-177;
parameter WEIGHT_0_193 = 16'd-2249;
parameter WEIGHT_0_194 = 16'd-1834;
parameter WEIGHT_0_195 = 16'd1763;
parameter WEIGHT_0_196 = 16'd458;
parameter WEIGHT_0_197 = 16'd-1355;
parameter WEIGHT_0_198 = 16'd489;
parameter WEIGHT_0_199 = 16'd2559;
parameter WEIGHT_0_200 = 16'd-2413;
parameter WEIGHT_0_201 = 16'd-1326;
parameter WEIGHT_0_202 = 16'd849;
parameter WEIGHT_0_203 = 16'd-1807;
parameter WEIGHT_0_204 = 16'd1512;
parameter WEIGHT_0_205 = 16'd-2564;
parameter WEIGHT_0_206 = 16'd-1962;
parameter WEIGHT_0_207 = 16'd2560;
parameter WEIGHT_0_208 = 16'd-500;
parameter WEIGHT_0_209 = 16'd2249;
parameter WEIGHT_0_210 = 16'd1788;
parameter WEIGHT_0_211 = 16'd-423;
parameter WEIGHT_0_212 = 16'd-1308;
parameter WEIGHT_0_213 = 16'd2143;
parameter WEIGHT_0_214 = 16'd-959;
parameter WEIGHT_0_215 = 16'd-1747;
parameter WEIGHT_0_216 = 16'd903;
parameter WEIGHT_0_217 = 16'd962;
parameter WEIGHT_0_218 = 16'd892;
parameter WEIGHT_0_219 = 16'd-538;
parameter WEIGHT_0_220 = 16'd-994;
parameter WEIGHT_0_221 = 16'd253;
parameter WEIGHT_0_222 = 16'd1547;
parameter WEIGHT_0_223 = 16'd672;
parameter WEIGHT_0_224 = 16'd2171;
parameter WEIGHT_0_225 = 16'd-2157;
parameter WEIGHT_0_226 = 16'd669;
parameter WEIGHT_0_227 = 16'd-1222;
parameter WEIGHT_0_228 = 16'd1767;
parameter WEIGHT_0_229 = 16'd561;
parameter WEIGHT_0_230 = 16'd-729;
parameter WEIGHT_0_231 = 16'd150;
parameter WEIGHT_0_232 = 16'd-2568;
parameter WEIGHT_0_233 = 16'd887;
parameter WEIGHT_0_234 = 16'd1234;
parameter WEIGHT_0_235 = 16'd1681;
parameter WEIGHT_0_236 = 16'd-251;
parameter WEIGHT_0_237 = 16'd-623;
parameter WEIGHT_0_238 = 16'd-2261;
parameter WEIGHT_0_239 = 16'd-1983;
parameter WEIGHT_0_240 = 16'd2006;
parameter WEIGHT_0_241 = 16'd658;
parameter WEIGHT_0_242 = 16'd2650;
parameter WEIGHT_0_243 = 16'd-2544;
parameter WEIGHT_0_244 = 16'd-2080;
parameter WEIGHT_0_245 = 16'd-133;
parameter WEIGHT_0_246 = 16'd570;
parameter WEIGHT_0_247 = 16'd-361;
parameter WEIGHT_0_248 = 16'd1337;
parameter WEIGHT_0_249 = 16'd-954;
parameter WEIGHT_0_250 = 16'd-1017;
parameter WEIGHT_0_251 = 16'd2140;
parameter WEIGHT_0_252 = 16'd144;
parameter WEIGHT_0_253 = 16'd-2090;
parameter WEIGHT_0_254 = 16'd2706;
parameter WEIGHT_0_255 = 16'd-1288;
parameter WEIGHT_0_256 = 16'd158;
parameter WEIGHT_0_257 = 16'd1201;
parameter WEIGHT_0_258 = 16'd-1251;
parameter WEIGHT_0_259 = 16'd1704;
parameter WEIGHT_0_260 = 16'd-1652;
parameter WEIGHT_0_261 = 16'd-167;
parameter WEIGHT_0_262 = 16'd-816;
parameter WEIGHT_0_263 = 16'd-439;
parameter WEIGHT_0_264 = 16'd-816;
parameter WEIGHT_0_265 = 16'd1302;
parameter WEIGHT_0_266 = 16'd11;
parameter WEIGHT_0_267 = 16'd1700;
parameter WEIGHT_0_268 = 16'd1420;
parameter WEIGHT_0_269 = 16'd-1764;
parameter WEIGHT_0_270 = 16'd2125;
parameter WEIGHT_0_271 = 16'd-1646;
parameter WEIGHT_0_272 = 16'd-1654;
parameter WEIGHT_0_273 = 16'd-2116;
parameter WEIGHT_0_274 = 16'd1352;
parameter WEIGHT_0_275 = 16'd-1165;
parameter WEIGHT_0_276 = 16'd-173;
parameter WEIGHT_0_277 = 16'd-2459;
parameter WEIGHT_0_278 = 16'd-1926;
parameter WEIGHT_0_279 = 16'd-84;
parameter WEIGHT_0_280 = 16'd1537;
parameter WEIGHT_0_281 = 16'd-1454;
parameter WEIGHT_0_282 = 16'd379;
parameter WEIGHT_0_283 = 16'd2054;
parameter WEIGHT_0_284 = 16'd1243;
parameter WEIGHT_0_285 = 16'd1484;
parameter WEIGHT_0_286 = 16'd-450;
parameter WEIGHT_0_287 = 16'd-522;
parameter WEIGHT_0_288 = 16'd-1299;
parameter WEIGHT_0_289 = 16'd276;
parameter WEIGHT_0_290 = 16'd1258;
parameter WEIGHT_0_291 = 16'd-2385;
parameter WEIGHT_0_292 = 16'd-2400;
parameter WEIGHT_0_293 = 16'd-1716;
parameter WEIGHT_0_294 = 16'd-1515;
parameter WEIGHT_0_295 = 16'd913;
parameter WEIGHT_0_296 = 16'd-1963;
parameter WEIGHT_0_297 = 16'd1190;
parameter WEIGHT_0_298 = 16'd2352;
parameter WEIGHT_0_299 = 16'd-1016;
parameter WEIGHT_0_300 = 16'd-1233;
parameter WEIGHT_0_301 = 16'd459;
parameter WEIGHT_0_302 = 16'd938;
parameter WEIGHT_0_303 = 16'd1869;
parameter WEIGHT_0_304 = 16'd-2061;
parameter WEIGHT_0_305 = 16'd-2790;
parameter WEIGHT_0_306 = 16'd-728;
parameter WEIGHT_0_307 = 16'd1276;
parameter WEIGHT_0_308 = 16'd-1391;
parameter WEIGHT_0_309 = 16'd-2281;
parameter WEIGHT_0_310 = 16'd-317;
parameter WEIGHT_0_311 = 16'd838;
parameter WEIGHT_0_312 = 16'd1747;
parameter WEIGHT_0_313 = 16'd-2569;
parameter WEIGHT_0_314 = 16'd-470;
parameter WEIGHT_0_315 = 16'd-1331;
parameter WEIGHT_0_316 = 16'd2791;
parameter WEIGHT_0_317 = 16'd1108;
parameter WEIGHT_0_318 = 16'd806;
parameter WEIGHT_0_319 = 16'd1160;
parameter WEIGHT_0_320 = 16'd180;
parameter WEIGHT_0_321 = 16'd-2451;
parameter WEIGHT_0_322 = 16'd-2214;
parameter WEIGHT_0_323 = 16'd-1775;
parameter WEIGHT_0_324 = 16'd-2780;
parameter WEIGHT_0_325 = 16'd-1023;
parameter WEIGHT_0_326 = 16'd176;
parameter WEIGHT_0_327 = 16'd2703;
parameter WEIGHT_0_328 = 16'd-2883;
parameter WEIGHT_0_329 = 16'd628;
parameter WEIGHT_0_330 = 16'd2470;
parameter WEIGHT_0_331 = 16'd1599;
parameter WEIGHT_0_332 = 16'd-3927;
parameter WEIGHT_0_333 = 16'd-708;
parameter WEIGHT_0_334 = 16'd-5065;
parameter WEIGHT_0_335 = 16'd620;
parameter WEIGHT_0_336 = 16'd1709;
parameter WEIGHT_0_337 = 16'd-1182;
parameter WEIGHT_0_338 = 16'd1489;
parameter WEIGHT_0_339 = 16'd1672;
parameter WEIGHT_0_340 = 16'd160;
parameter WEIGHT_0_341 = 16'd1215;
parameter WEIGHT_0_342 = 16'd-3761;
parameter WEIGHT_0_343 = 16'd-1380;
parameter WEIGHT_0_344 = 16'd-4612;
parameter WEIGHT_0_345 = 16'd-558;
parameter WEIGHT_0_346 = 16'd5875;
parameter WEIGHT_0_347 = 16'd959;
parameter WEIGHT_0_348 = 16'd-2243;
parameter WEIGHT_0_349 = 16'd1399;
parameter WEIGHT_0_350 = 16'd1938;
parameter WEIGHT_0_351 = 16'd1511;
parameter WEIGHT_0_352 = 16'd-4062;
parameter WEIGHT_0_353 = 16'd423;
parameter WEIGHT_0_354 = 16'd-6968;
parameter WEIGHT_0_355 = 16'd-2846;
parameter WEIGHT_0_356 = 16'd2888;
parameter WEIGHT_0_357 = 16'd-152;
parameter WEIGHT_0_358 = 16'd1623;
parameter WEIGHT_0_359 = 16'd-505;
parameter WEIGHT_0_360 = 16'd-376;
parameter WEIGHT_0_361 = 16'd-4798;
parameter WEIGHT_0_362 = 16'd-4112;
parameter WEIGHT_0_363 = 16'd-4341;
parameter WEIGHT_0_364 = 16'd-6086;
parameter WEIGHT_0_365 = 16'd-1812;
parameter WEIGHT_0_366 = 16'd5521;
parameter WEIGHT_0_367 = 16'd-773;
parameter WEIGHT_0_368 = 16'd-4081;
parameter WEIGHT_0_369 = 16'd-6863;
parameter WEIGHT_0_370 = 16'd-1474;
parameter WEIGHT_0_371 = 16'd-1427;
parameter WEIGHT_0_372 = 16'd-2473;
parameter WEIGHT_0_373 = 16'd-1533;
parameter WEIGHT_0_374 = 16'd-8403;
parameter WEIGHT_0_375 = 16'd-3287;
parameter WEIGHT_0_376 = 16'd6445;
parameter WEIGHT_0_377 = 16'd-5297;
parameter WEIGHT_0_378 = 16'd-4024;
parameter WEIGHT_0_379 = 16'd-4325;
parameter WEIGHT_0_380 = 16'd-970;
parameter WEIGHT_0_381 = 16'd-2458;
parameter WEIGHT_0_382 = 16'd-5622;
parameter WEIGHT_0_383 = 16'd-1977;
parameter WEIGHT_0_384 = 16'd-8395;
parameter WEIGHT_0_385 = 16'd-540;
parameter WEIGHT_0_386 = 16'd4310;
parameter WEIGHT_0_387 = 16'd-4884;
parameter WEIGHT_0_388 = 16'd-972;
parameter WEIGHT_0_389 = 16'd-3115;
parameter WEIGHT_0_390 = 16'd-1347;
parameter WEIGHT_0_391 = 16'd-4380;
parameter WEIGHT_0_392 = 16'd-7898;
parameter WEIGHT_0_393 = 16'd-3839;
parameter WEIGHT_0_394 = 16'd-10564;
parameter WEIGHT_0_395 = 16'd-3739;
parameter WEIGHT_0_396 = 16'd10895;
parameter WEIGHT_0_397 = 16'd-6181;
parameter WEIGHT_0_398 = 16'd-7708;
parameter WEIGHT_0_399 = 16'd-8296;
parameter WEIGHT_0_400 = 16'd2553;
parameter WEIGHT_0_401 = 16'd-3558;
parameter WEIGHT_0_402 = 16'd-8723;
parameter WEIGHT_0_403 = 16'd-3687;
parameter WEIGHT_0_404 = 16'd-13983;
parameter WEIGHT_0_405 = 16'd-2781;
parameter WEIGHT_0_406 = 16'd7706;
parameter WEIGHT_0_407 = 16'd-7190;
parameter WEIGHT_0_408 = 16'd-6234;
parameter WEIGHT_0_409 = 16'd-9164;
parameter WEIGHT_0_410 = 16'd2141;
parameter WEIGHT_0_411 = 16'd-3510;
parameter WEIGHT_0_412 = 16'd-5501;
parameter WEIGHT_0_413 = 16'd-2962;
parameter WEIGHT_0_414 = 16'd-12023;
parameter WEIGHT_0_415 = 16'd-4349;
parameter WEIGHT_0_416 = 16'd10238;
parameter WEIGHT_0_417 = 16'd-1176;
parameter WEIGHT_0_418 = 16'd-4853;
parameter WEIGHT_0_419 = 16'd-5763;
parameter WEIGHT_0_420 = 16'd-4097;
parameter WEIGHT_0_421 = 16'd4422;
parameter WEIGHT_0_422 = 16'd-1273;
parameter WEIGHT_0_423 = 16'd-4631;
parameter WEIGHT_0_424 = 16'd-3587;
parameter WEIGHT_0_425 = 16'd-3235;
parameter WEIGHT_0_426 = 16'd-717;
parameter WEIGHT_0_427 = 16'd-3477;
parameter WEIGHT_0_428 = 16'd-5401;
parameter WEIGHT_0_429 = 16'd-5673;
parameter WEIGHT_0_430 = 16'd2783;
parameter WEIGHT_0_431 = 16'd-403;
parameter WEIGHT_0_432 = 16'd393;
parameter WEIGHT_0_433 = 16'd-2116;
parameter WEIGHT_0_434 = 16'd-10246;
parameter WEIGHT_0_435 = 16'd-6343;
parameter WEIGHT_0_436 = 16'd2005;
parameter WEIGHT_0_437 = 16'd-2630;
parameter WEIGHT_0_438 = 16'd-1534;
parameter WEIGHT_0_439 = 16'd-7638;
parameter WEIGHT_0_440 = 16'd-1382;
parameter WEIGHT_0_441 = 16'd-5055;
parameter WEIGHT_0_442 = 16'd6632;
parameter WEIGHT_0_443 = 16'd-5702;
parameter WEIGHT_0_444 = 16'd-14503;
parameter WEIGHT_0_445 = 16'd-10282;
parameter WEIGHT_0_446 = 16'd1222;
parameter WEIGHT_0_447 = 16'd-4500;
parameter WEIGHT_0_448 = 16'd-8018;
parameter WEIGHT_0_449 = 16'd-5326;
parameter WEIGHT_0_450 = 16'd680;
parameter WEIGHT_0_451 = 16'd-7004;
parameter WEIGHT_0_452 = 16'd2959;
parameter WEIGHT_0_453 = 16'd-2492;
parameter WEIGHT_0_454 = 16'd-9423;
parameter WEIGHT_0_455 = 16'd-3151;
parameter WEIGHT_0_456 = 16'd3734;
parameter WEIGHT_0_457 = 16'd-192;
parameter WEIGHT_0_458 = 16'd-6732;
parameter WEIGHT_0_459 = 16'd-5417;
parameter WEIGHT_0_460 = 16'd-3859;
parameter WEIGHT_0_461 = 16'd595;
parameter WEIGHT_0_462 = 16'd-6214;
parameter WEIGHT_0_463 = 16'd-460;
parameter WEIGHT_0_464 = 16'd-9320;
parameter WEIGHT_0_465 = 16'd-2917;
parameter WEIGHT_0_466 = 16'd7970;
parameter WEIGHT_0_467 = 16'd-876;
parameter WEIGHT_0_468 = 16'd-1937;
parameter WEIGHT_0_469 = 16'd-3949;
parameter WEIGHT_0_470 = 16'd-4849;
parameter WEIGHT_0_471 = 16'd-459;
parameter WEIGHT_0_472 = 16'd-9106;
parameter WEIGHT_0_473 = 16'd-896;
parameter WEIGHT_0_474 = 16'd-9870;
parameter WEIGHT_0_475 = 16'd-9771;
parameter WEIGHT_0_476 = 16'd7927;
parameter WEIGHT_0_477 = 16'd-6598;
parameter WEIGHT_0_478 = 16'd-8366;
parameter WEIGHT_0_479 = 16'd-9080;
parameter WEIGHT_0_480 = 16'd-860;
parameter WEIGHT_0_481 = 16'd-3191;
parameter WEIGHT_0_482 = 16'd-8581;
parameter WEIGHT_0_483 = 16'd-205;
parameter WEIGHT_0_484 = 16'd-10185;
parameter WEIGHT_0_485 = 16'd-4675;
parameter WEIGHT_0_486 = 16'd6988;
parameter WEIGHT_0_487 = 16'd-2818;
parameter WEIGHT_0_488 = 16'd-4114;
parameter WEIGHT_0_489 = 16'd-8559;
parameter WEIGHT_0_490 = 16'd-1630;
parameter WEIGHT_0_491 = 16'd504;
parameter WEIGHT_0_492 = 16'd-6126;
parameter WEIGHT_0_493 = 16'd-2519;
parameter WEIGHT_0_494 = 16'd-3605;
parameter WEIGHT_0_495 = 16'd-4123;
parameter WEIGHT_0_496 = 16'd5455;
parameter WEIGHT_0_497 = 16'd144;
parameter WEIGHT_0_498 = 16'd-4481;
parameter WEIGHT_0_499 = 16'd-5481;
parameter WEIGHT_0_500 = 16'd-3393;
parameter WEIGHT_0_501 = 16'd540;
parameter WEIGHT_0_502 = 16'd-4886;
parameter WEIGHT_0_503 = 16'd589;
parameter WEIGHT_0_504 = 16'd-2372;
parameter WEIGHT_0_505 = 16'd-1577;
parameter WEIGHT_0_506 = 16'd3596;
parameter WEIGHT_0_507 = 16'd-2259;
parameter WEIGHT_0_508 = 16'd-5006;
parameter WEIGHT_0_509 = 16'd-4807;
parameter WEIGHT_0_510 = 16'd-1089;
parameter WEIGHT_0_511 = 16'd-2493;
parameter WEIGHT_0_512 = 16'd-1675;
parameter WEIGHT_0_513 = 16'd-163;
parameter WEIGHT_0_514 = 16'd-3763;
parameter WEIGHT_0_515 = 16'd-1796;
parameter WEIGHT_0_516 = 16'd3234;
parameter WEIGHT_0_517 = 16'd-3440;
parameter WEIGHT_0_518 = 16'd-3022;
parameter WEIGHT_0_519 = 16'd-3142;
parameter WEIGHT_0_520 = 16'd-1092;
parameter WEIGHT_0_521 = 16'd2668;
parameter WEIGHT_0_522 = 16'd2218;
parameter WEIGHT_0_523 = 16'd-2579;
parameter WEIGHT_0_524 = 16'd-1828;
parameter WEIGHT_0_525 = 16'd-1224;
parameter WEIGHT_0_526 = 16'd-965;
parameter WEIGHT_0_527 = 16'd-2428;
parameter WEIGHT_0_528 = 16'd-472;
parameter WEIGHT_0_529 = 16'd-254;
parameter WEIGHT_0_530 = 16'd-1200;
parameter WEIGHT_0_531 = 16'd370;
parameter WEIGHT_0_532 = 16'd2242;
parameter WEIGHT_0_533 = 16'd2169;
parameter WEIGHT_0_534 = 16'd2798;
parameter WEIGHT_0_535 = 16'd-1304;
parameter WEIGHT_0_536 = 16'd-24;
parameter WEIGHT_0_537 = 16'd585;
parameter WEIGHT_0_538 = 16'd-2393;
parameter WEIGHT_0_539 = 16'd-2603;
parameter WEIGHT_0_540 = 16'd2107;
parameter WEIGHT_0_541 = 16'd2077;
parameter WEIGHT_0_542 = 16'd755;
parameter WEIGHT_0_543 = 16'd2339;
parameter WEIGHT_0_544 = 16'd-491;
parameter WEIGHT_0_545 = 16'd-2624;
parameter WEIGHT_0_546 = 16'd1310;
parameter WEIGHT_0_547 = 16'd2761;
parameter WEIGHT_0_548 = 16'd2048;
parameter WEIGHT_0_549 = 16'd985;
parameter WEIGHT_0_550 = 16'd-2090;
parameter WEIGHT_0_551 = 16'd773;
parameter WEIGHT_0_552 = 16'd425;
parameter WEIGHT_0_553 = 16'd-1506;
parameter WEIGHT_0_554 = 16'd-410;
parameter WEIGHT_0_555 = 16'd-1596;
parameter WEIGHT_0_556 = 16'd2108;
parameter WEIGHT_0_557 = 16'd-15;
parameter WEIGHT_0_558 = 16'd605;
parameter WEIGHT_0_559 = 16'd-2023;
parameter WEIGHT_0_560 = 16'd-2652;
parameter WEIGHT_0_561 = 16'd-837;
parameter WEIGHT_0_562 = 16'd-141;
parameter WEIGHT_0_563 = 16'd2012;
parameter WEIGHT_0_564 = 16'd225;
parameter WEIGHT_0_565 = 16'd-913;
parameter WEIGHT_0_566 = 16'd1451;
parameter WEIGHT_0_567 = 16'd-1089;
parameter WEIGHT_0_568 = 16'd-2337;
parameter WEIGHT_0_569 = 16'd-1689;
parameter WEIGHT_0_570 = 16'd-2543;
parameter WEIGHT_0_571 = 16'd375;
parameter WEIGHT_0_572 = 16'd2533;
parameter WEIGHT_0_573 = 16'd-411;
parameter WEIGHT_0_574 = 16'd-1044;
parameter WEIGHT_0_575 = 16'd-108;
parameter WEIGHT_0_576 = 16'd-2033;
parameter WEIGHT_0_577 = 16'd455;
parameter WEIGHT_0_578 = 16'd981;
parameter WEIGHT_0_579 = 16'd2692;
parameter WEIGHT_0_580 = 16'd2049;
parameter WEIGHT_0_581 = 16'd-1205;
parameter WEIGHT_0_582 = 16'd133;
parameter WEIGHT_0_583 = 16'd-1895;
parameter WEIGHT_0_584 = 16'd-2381;
parameter WEIGHT_0_585 = 16'd-1755;
parameter WEIGHT_0_586 = 16'd272;
parameter WEIGHT_0_587 = 16'd-2777;
parameter WEIGHT_0_588 = 16'd1995;
parameter WEIGHT_0_589 = 16'd-600;
parameter WEIGHT_0_590 = 16'd1688;
parameter WEIGHT_0_591 = 16'd-1323;
parameter WEIGHT_0_592 = 16'd-3382;
parameter WEIGHT_0_593 = 16'd-3559;
parameter WEIGHT_0_594 = 16'd-4304;
parameter WEIGHT_0_595 = 16'd-4103;
parameter WEIGHT_0_596 = 16'd2225;
parameter WEIGHT_0_597 = 16'd-2898;
parameter WEIGHT_0_598 = 16'd-1748;
parameter WEIGHT_0_599 = 16'd476;
parameter WEIGHT_0_600 = 16'd-238;
parameter WEIGHT_0_601 = 16'd1082;
parameter WEIGHT_0_602 = 16'd-2062;
parameter WEIGHT_0_603 = 16'd-424;
parameter WEIGHT_0_604 = 16'd-7195;
parameter WEIGHT_0_605 = 16'd-3995;
parameter WEIGHT_0_606 = 16'd2662;
parameter WEIGHT_0_607 = 16'd-2940;
parameter WEIGHT_0_608 = 16'd-2590;
parameter WEIGHT_0_609 = 16'd50;
parameter WEIGHT_0_610 = 16'd-4188;
parameter WEIGHT_0_611 = 16'd-1909;
parameter WEIGHT_0_612 = 16'd-3325;
parameter WEIGHT_0_613 = 16'd-998;
parameter WEIGHT_0_614 = 16'd-155;
parameter WEIGHT_0_615 = 16'd661;
parameter WEIGHT_0_616 = 16'd1277;
parameter WEIGHT_0_617 = 16'd-1963;
parameter WEIGHT_0_618 = 16'd-572;
parameter WEIGHT_0_619 = 16'd1138;
parameter WEIGHT_0_620 = 16'd-5069;
parameter WEIGHT_0_621 = 16'd587;
parameter WEIGHT_0_622 = 16'd-834;
parameter WEIGHT_0_623 = 16'd-949;
parameter WEIGHT_0_624 = 16'd-7850;
parameter WEIGHT_0_625 = 16'd837;
parameter WEIGHT_0_626 = 16'd5908;
parameter WEIGHT_0_627 = 16'd1618;
parameter WEIGHT_0_628 = 16'd1019;
parameter WEIGHT_0_629 = 16'd-277;
parameter WEIGHT_0_630 = 16'd-6082;
parameter WEIGHT_0_631 = 16'd-2249;
parameter WEIGHT_0_632 = 16'd-2672;
parameter WEIGHT_0_633 = 16'd-2658;
parameter WEIGHT_0_634 = 16'd-9450;
parameter WEIGHT_0_635 = 16'd-1033;
parameter WEIGHT_0_636 = 16'd6784;
parameter WEIGHT_0_637 = 16'd-2576;
parameter WEIGHT_0_638 = 16'd-6796;
parameter WEIGHT_0_639 = 16'd-1960;
parameter WEIGHT_0_640 = 16'd-4769;
parameter WEIGHT_0_641 = 16'd-7174;
parameter WEIGHT_0_642 = 16'd-621;
parameter WEIGHT_0_643 = 16'd-5500;
parameter WEIGHT_0_644 = 16'd-14708;
parameter WEIGHT_0_645 = 16'd-7450;
parameter WEIGHT_0_646 = 16'd9407;
parameter WEIGHT_0_647 = 16'd-6891;
parameter WEIGHT_0_648 = 16'd-9623;
parameter WEIGHT_0_649 = 16'd-5549;
parameter WEIGHT_0_650 = 16'd-11961;
parameter WEIGHT_0_651 = 16'd-4453;
parameter WEIGHT_0_652 = 16'd-214;
parameter WEIGHT_0_653 = 16'd-11553;
parameter WEIGHT_0_654 = 16'd-18390;
parameter WEIGHT_0_655 = 16'd-5624;
parameter WEIGHT_0_656 = 16'd7460;
parameter WEIGHT_0_657 = 16'd-8402;
parameter WEIGHT_0_658 = 16'd-8551;
parameter WEIGHT_0_659 = 16'd-7086;
parameter WEIGHT_0_660 = 16'd-10963;
parameter WEIGHT_0_661 = 16'd-7993;
parameter WEIGHT_0_662 = 16'd2115;
parameter WEIGHT_0_663 = 16'd-4268;
parameter WEIGHT_0_664 = 16'd-18696;
parameter WEIGHT_0_665 = 16'd-7459;
parameter WEIGHT_0_666 = 16'd8831;
parameter WEIGHT_0_667 = 16'd-8551;
parameter WEIGHT_0_668 = 16'd-14727;
parameter WEIGHT_0_669 = 16'd-12683;
parameter WEIGHT_0_670 = 16'd-6629;
parameter WEIGHT_0_671 = 16'd-7261;
parameter WEIGHT_0_672 = 16'd210;
parameter WEIGHT_0_673 = 16'd221;
parameter WEIGHT_0_674 = 16'd-22592;
parameter WEIGHT_0_675 = 16'd-7094;
parameter WEIGHT_0_676 = 16'd13435;
parameter WEIGHT_0_677 = 16'd-7626;
parameter WEIGHT_0_678 = 16'd-20656;
parameter WEIGHT_0_679 = 16'd-16800;
parameter WEIGHT_0_680 = 16'd-8435;
parameter WEIGHT_0_681 = 16'd-2291;
parameter WEIGHT_0_682 = 16'd1839;
parameter WEIGHT_0_683 = 16'd-167;
parameter WEIGHT_0_684 = 16'd-20747;
parameter WEIGHT_0_685 = 16'd-11606;
parameter WEIGHT_0_686 = 16'd11163;
parameter WEIGHT_0_687 = 16'd-9816;
parameter WEIGHT_0_688 = 16'd-18560;
parameter WEIGHT_0_689 = 16'd-14089;
parameter WEIGHT_0_690 = 16'd-9652;
parameter WEIGHT_0_691 = 16'd3904;
parameter WEIGHT_0_692 = 16'd1711;
parameter WEIGHT_0_693 = 16'd-3097;
parameter WEIGHT_0_694 = 16'd-16843;
parameter WEIGHT_0_695 = 16'd-16668;
parameter WEIGHT_0_696 = 16'd7857;
parameter WEIGHT_0_697 = 16'd-11297;
parameter WEIGHT_0_698 = 16'd-20543;
parameter WEIGHT_0_699 = 16'd-18023;
parameter WEIGHT_0_700 = 16'd-12024;
parameter WEIGHT_0_701 = 16'd1552;
parameter WEIGHT_0_702 = 16'd310;
parameter WEIGHT_0_703 = 16'd-4514;
parameter WEIGHT_0_704 = 16'd-13139;
parameter WEIGHT_0_705 = 16'd-17298;
parameter WEIGHT_0_706 = 16'd8039;
parameter WEIGHT_0_707 = 16'd-5235;
parameter WEIGHT_0_708 = 16'd-21917;
parameter WEIGHT_0_709 = 16'd-13470;
parameter WEIGHT_0_710 = 16'd-16567;
parameter WEIGHT_0_711 = 16'd4262;
parameter WEIGHT_0_712 = 16'd1648;
parameter WEIGHT_0_713 = 16'd-6582;
parameter WEIGHT_0_714 = 16'd-12885;
parameter WEIGHT_0_715 = 16'd-10613;
parameter WEIGHT_0_716 = 16'd4780;
parameter WEIGHT_0_717 = 16'd-6050;
parameter WEIGHT_0_718 = 16'd-17421;
parameter WEIGHT_0_719 = 16'd-16427;
parameter WEIGHT_0_720 = 16'd-13696;
parameter WEIGHT_0_721 = 16'd5280;
parameter WEIGHT_0_722 = 16'd2911;
parameter WEIGHT_0_723 = 16'd-5901;
parameter WEIGHT_0_724 = 16'd-15264;
parameter WEIGHT_0_725 = 16'd-5676;
parameter WEIGHT_0_726 = 16'd3705;
parameter WEIGHT_0_727 = 16'd-5108;
parameter WEIGHT_0_728 = 16'd-24737;
parameter WEIGHT_0_729 = 16'd-13447;
parameter WEIGHT_0_730 = 16'd-17873;
parameter WEIGHT_0_731 = 16'd-2990;
parameter WEIGHT_0_732 = 16'd2995;
parameter WEIGHT_0_733 = 16'd-6769;
parameter WEIGHT_0_734 = 16'd-10035;
parameter WEIGHT_0_735 = 16'd1087;
parameter WEIGHT_0_736 = 16'd6452;
parameter WEIGHT_0_737 = 16'd-6468;
parameter WEIGHT_0_738 = 16'd-14837;
parameter WEIGHT_0_739 = 16'd-9780;
parameter WEIGHT_0_740 = 16'd-16793;
parameter WEIGHT_0_741 = 16'd-4301;
parameter WEIGHT_0_742 = 16'd-2126;
parameter WEIGHT_0_743 = 16'd-5829;
parameter WEIGHT_0_744 = 16'd-21359;
parameter WEIGHT_0_745 = 16'd-394;
parameter WEIGHT_0_746 = 16'd6741;
parameter WEIGHT_0_747 = 16'd-1628;
parameter WEIGHT_0_748 = 16'd-6381;
parameter WEIGHT_0_749 = 16'd-7882;
parameter WEIGHT_0_750 = 16'd-13612;
parameter WEIGHT_0_751 = 16'd-1110;
parameter WEIGHT_0_752 = 16'd-9237;
parameter WEIGHT_0_753 = 16'd-6294;
parameter WEIGHT_0_754 = 16'd-9418;
parameter WEIGHT_0_755 = 16'd-545;
parameter WEIGHT_0_756 = 16'd7600;
parameter WEIGHT_0_757 = 16'd-3982;
parameter WEIGHT_0_758 = 16'd-16429;
parameter WEIGHT_0_759 = 16'd-11046;
parameter WEIGHT_0_760 = 16'd-15793;
parameter WEIGHT_0_761 = 16'd-3479;
parameter WEIGHT_0_762 = 16'd-4338;
parameter WEIGHT_0_763 = 16'd-5475;
parameter WEIGHT_0_764 = 16'd-6122;
parameter WEIGHT_0_765 = 16'd-5834;
parameter WEIGHT_0_766 = 16'd7155;
parameter WEIGHT_0_767 = 16'd-1960;
parameter WEIGHT_0_768 = 16'd-8324;
parameter WEIGHT_0_769 = 16'd-7805;
parameter WEIGHT_0_770 = 16'd-6708;
parameter WEIGHT_0_771 = 16'd-8309;
parameter WEIGHT_0_772 = 16'd-6089;
parameter WEIGHT_0_773 = 16'd-8103;
parameter WEIGHT_0_774 = 16'd-6185;
parameter WEIGHT_0_775 = 16'd-7194;
parameter WEIGHT_0_776 = 16'd7043;
parameter WEIGHT_0_777 = 16'd332;
parameter WEIGHT_0_778 = 16'd-8310;
parameter WEIGHT_0_779 = 16'd-3580;
parameter WEIGHT_0_780 = 16'd-8746;
parameter WEIGHT_0_781 = 16'd-4071;
parameter WEIGHT_0_782 = 16'd-8861;
parameter WEIGHT_0_783 = 16'd-9965;
parameter WEIGHT_0_784 = 16'd-7927;
parameter WEIGHT_0_785 = 16'd-2934;
parameter WEIGHT_0_786 = 16'd8236;
parameter WEIGHT_0_787 = 16'd-3970;
parameter WEIGHT_0_788 = 16'd-4616;
parameter WEIGHT_0_789 = 16'd-6323;
parameter WEIGHT_0_790 = 16'd-5408;
parameter WEIGHT_0_791 = 16'd-3656;
parameter WEIGHT_0_792 = 16'd-1539;
parameter WEIGHT_0_793 = 16'd-1960;
parameter WEIGHT_0_794 = 16'd-10040;
parameter WEIGHT_0_795 = 16'd-2955;
parameter WEIGHT_0_796 = 16'd8574;
parameter WEIGHT_0_797 = 16'd-536;
parameter WEIGHT_0_798 = 16'd-9237;
parameter WEIGHT_0_799 = 16'd-4238;
parameter WEIGHT_0_800 = 16'd-1091;
parameter WEIGHT_0_801 = 16'd-2299;
parameter WEIGHT_0_802 = 16'd4406;
parameter WEIGHT_0_803 = 16'd-2082;
parameter WEIGHT_0_804 = 16'd-7233;
parameter WEIGHT_0_805 = 16'd-7953;
parameter WEIGHT_0_806 = 16'd-2214;
parameter WEIGHT_0_807 = 16'd-1693;
parameter WEIGHT_0_808 = 16'd-2628;
parameter WEIGHT_0_809 = 16'd-203;
parameter WEIGHT_0_810 = 16'd-3858;
parameter WEIGHT_0_811 = 16'd-3129;
parameter WEIGHT_0_812 = 16'd-68;
parameter WEIGHT_0_813 = 16'd-1974;
parameter WEIGHT_0_814 = 16'd-3769;
parameter WEIGHT_0_815 = 16'd-3775;
parameter WEIGHT_0_816 = 16'd-2051;
parameter WEIGHT_0_817 = 16'd-2163;
parameter WEIGHT_0_818 = 16'd-4322;
parameter WEIGHT_0_819 = 16'd-2248;
parameter WEIGHT_0_820 = 16'd1226;
parameter WEIGHT_0_821 = 16'd-2044;
parameter WEIGHT_0_822 = 16'd-1908;
parameter WEIGHT_0_823 = 16'd-1046;
parameter WEIGHT_0_824 = 16'd2019;
parameter WEIGHT_0_825 = 16'd2717;
parameter WEIGHT_0_826 = 16'd2571;
parameter WEIGHT_0_827 = 16'd1784;
parameter WEIGHT_0_828 = 16'd-2379;
parameter WEIGHT_0_829 = 16'd-2758;
parameter WEIGHT_0_830 = 16'd-1083;
parameter WEIGHT_0_831 = 16'd-943;
parameter WEIGHT_0_832 = 16'd739;
parameter WEIGHT_0_833 = 16'd209;
parameter WEIGHT_0_834 = 16'd1239;
parameter WEIGHT_0_835 = 16'd548;
parameter WEIGHT_0_836 = 16'd512;
parameter WEIGHT_0_837 = 16'd-2672;
parameter WEIGHT_0_838 = 16'd1939;
parameter WEIGHT_0_839 = 16'd1097;
parameter WEIGHT_0_840 = 16'd1779;
parameter WEIGHT_0_841 = 16'd1543;
parameter WEIGHT_0_842 = 16'd2483;
parameter WEIGHT_0_843 = 16'd-16;
parameter WEIGHT_0_844 = 16'd-1816;
parameter WEIGHT_0_845 = 16'd2331;
parameter WEIGHT_0_846 = 16'd-831;
parameter WEIGHT_0_847 = 16'd-2169;
parameter WEIGHT_0_848 = 16'd-1547;
parameter WEIGHT_0_849 = 16'd-2271;
parameter WEIGHT_0_850 = 16'd2711;
parameter WEIGHT_0_851 = 16'd779;
parameter WEIGHT_0_852 = 16'd-1192;
parameter WEIGHT_0_853 = 16'd2199;
parameter WEIGHT_0_854 = 16'd-2685;
parameter WEIGHT_0_855 = 16'd1597;
parameter WEIGHT_0_856 = 16'd-1941;
parameter WEIGHT_0_857 = 16'd1482;
parameter WEIGHT_0_858 = 16'd-747;
parameter WEIGHT_0_859 = 16'd-2260;
parameter WEIGHT_0_860 = 16'd-220;
parameter WEIGHT_0_861 = 16'd3782;
parameter WEIGHT_0_862 = 16'd-3913;
parameter WEIGHT_0_863 = 16'd-689;
parameter WEIGHT_0_864 = 16'd-536;
parameter WEIGHT_0_865 = 16'd497;
parameter WEIGHT_0_866 = 16'd-360;
parameter WEIGHT_0_867 = 16'd1941;
parameter WEIGHT_0_868 = 16'd-4369;
parameter WEIGHT_0_869 = 16'd-1326;
parameter WEIGHT_0_870 = 16'd-758;
parameter WEIGHT_0_871 = 16'd599;
parameter WEIGHT_0_872 = 16'd-2580;
parameter WEIGHT_0_873 = 16'd-1465;
parameter WEIGHT_0_874 = 16'd-4210;
parameter WEIGHT_0_875 = 16'd-3050;
parameter WEIGHT_0_876 = 16'd1049;
parameter WEIGHT_0_877 = 16'd-492;
parameter WEIGHT_0_878 = 16'd-5420;
parameter WEIGHT_0_879 = 16'd-2707;
parameter WEIGHT_0_880 = 16'd-5932;
parameter WEIGHT_0_881 = 16'd-1738;
parameter WEIGHT_0_882 = 16'd-6132;
parameter WEIGHT_0_883 = 16'd-6033;
parameter WEIGHT_0_884 = 16'd-5536;
parameter WEIGHT_0_885 = 16'd1628;
parameter WEIGHT_0_886 = 16'd4606;
parameter WEIGHT_0_887 = 16'd-5300;
parameter WEIGHT_0_888 = 16'd-5102;
parameter WEIGHT_0_889 = 16'd-5384;
parameter WEIGHT_0_890 = 16'd-1888;
parameter WEIGHT_0_891 = 16'd-3007;
parameter WEIGHT_0_892 = 16'd-3746;
parameter WEIGHT_0_893 = 16'd5279;
parameter WEIGHT_0_894 = 16'd-3388;
parameter WEIGHT_0_895 = 16'd-3041;
parameter WEIGHT_0_896 = 16'd5740;
parameter WEIGHT_0_897 = 16'd-4820;
parameter WEIGHT_0_898 = 16'd-10583;
parameter WEIGHT_0_899 = 16'd-4882;
parameter WEIGHT_0_900 = 16'd-4448;
parameter WEIGHT_0_901 = 16'd-5225;
parameter WEIGHT_0_902 = 16'd3000;
parameter WEIGHT_0_903 = 16'd3725;
parameter WEIGHT_0_904 = 16'd-6385;
parameter WEIGHT_0_905 = 16'd-3534;
parameter WEIGHT_0_906 = 16'd7300;
parameter WEIGHT_0_907 = 16'd-5598;
parameter WEIGHT_0_908 = 16'd-4907;
parameter WEIGHT_0_909 = 16'd-755;
parameter WEIGHT_0_910 = 16'd-8460;
parameter WEIGHT_0_911 = 16'd-5405;
parameter WEIGHT_0_912 = 16'd2920;
parameter WEIGHT_0_913 = 16'd4633;
parameter WEIGHT_0_914 = 16'd-9800;
parameter WEIGHT_0_915 = 16'd-9195;
parameter WEIGHT_0_916 = 16'd8396;
parameter WEIGHT_0_917 = 16'd-8048;
parameter WEIGHT_0_918 = 16'd-7945;
parameter WEIGHT_0_919 = 16'd-6053;
parameter WEIGHT_0_920 = 16'd-6786;
parameter WEIGHT_0_921 = 16'd-12802;
parameter WEIGHT_0_922 = 16'd3128;
parameter WEIGHT_0_923 = 16'd1317;
parameter WEIGHT_0_924 = 16'd-11674;
parameter WEIGHT_0_925 = 16'd-7062;
parameter WEIGHT_0_926 = 16'd4275;
parameter WEIGHT_0_927 = 16'd-11530;
parameter WEIGHT_0_928 = 16'd-6175;
parameter WEIGHT_0_929 = 16'd-10826;
parameter WEIGHT_0_930 = 16'd-4642;
parameter WEIGHT_0_931 = 16'd-9207;
parameter WEIGHT_0_932 = 16'd8848;
parameter WEIGHT_0_933 = 16'd-773;
parameter WEIGHT_0_934 = 16'd-15080;
parameter WEIGHT_0_935 = 16'd-5996;
parameter WEIGHT_0_936 = 16'd6878;
parameter WEIGHT_0_937 = 16'd-14466;
parameter WEIGHT_0_938 = 16'd-11370;
parameter WEIGHT_0_939 = 16'd-10272;
parameter WEIGHT_0_940 = 16'd-6659;
parameter WEIGHT_0_941 = 16'd-12753;
parameter WEIGHT_0_942 = 16'd5559;
parameter WEIGHT_0_943 = 16'd2582;
parameter WEIGHT_0_944 = 16'd-18176;
parameter WEIGHT_0_945 = 16'd-5317;
parameter WEIGHT_0_946 = 16'd7410;
parameter WEIGHT_0_947 = 16'd-16164;
parameter WEIGHT_0_948 = 16'd-13135;
parameter WEIGHT_0_949 = 16'd-15681;
parameter WEIGHT_0_950 = 16'd-3409;
parameter WEIGHT_0_951 = 16'd-15182;
parameter WEIGHT_0_952 = 16'd7747;
parameter WEIGHT_0_953 = 16'd6838;
parameter WEIGHT_0_954 = 16'd-23785;
parameter WEIGHT_0_955 = 16'd-6283;
parameter WEIGHT_0_956 = 16'd5493;
parameter WEIGHT_0_957 = 16'd-17568;
parameter WEIGHT_0_958 = 16'd-9547;
parameter WEIGHT_0_959 = 16'd-18919;
parameter WEIGHT_0_960 = 16'd-5692;
parameter WEIGHT_0_961 = 16'd-10686;
parameter WEIGHT_0_962 = 16'd9301;
parameter WEIGHT_0_963 = 16'd10002;
parameter WEIGHT_0_964 = 16'd-25743;
parameter WEIGHT_0_965 = 16'd-6212;
parameter WEIGHT_0_966 = 16'd2374;
parameter WEIGHT_0_967 = 16'd-16912;
parameter WEIGHT_0_968 = 16'd-13596;
parameter WEIGHT_0_969 = 16'd-20365;
parameter WEIGHT_0_970 = 16'd-915;
parameter WEIGHT_0_971 = 16'd-2895;
parameter WEIGHT_0_972 = 16'd9235;
parameter WEIGHT_0_973 = 16'd8315;
parameter WEIGHT_0_974 = 16'd-23098;
parameter WEIGHT_0_975 = 16'd-3455;
parameter WEIGHT_0_976 = 16'd7840;
parameter WEIGHT_0_977 = 16'd-17496;
parameter WEIGHT_0_978 = 16'd-6586;
parameter WEIGHT_0_979 = 16'd-24264;
parameter WEIGHT_0_980 = 16'd-3756;
parameter WEIGHT_0_981 = 16'd-4067;
parameter WEIGHT_0_982 = 16'd6179;
parameter WEIGHT_0_983 = 16'd6691;
parameter WEIGHT_0_984 = 16'd-16104;
parameter WEIGHT_0_985 = 16'd-2981;
parameter WEIGHT_0_986 = 16'd5408;
parameter WEIGHT_0_987 = 16'd-14309;
parameter WEIGHT_0_988 = 16'd-8212;
parameter WEIGHT_0_989 = 16'd-28387;
parameter WEIGHT_0_990 = 16'd-3886;
parameter WEIGHT_0_991 = 16'd-110;
parameter WEIGHT_0_992 = 16'd2790;
parameter WEIGHT_0_993 = 16'd5313;
parameter WEIGHT_0_994 = 16'd-16716;
parameter WEIGHT_0_995 = 16'd-412;
parameter WEIGHT_0_996 = 16'd4407;
parameter WEIGHT_0_997 = 16'd-15224;
parameter WEIGHT_0_998 = 16'd-10223;
parameter WEIGHT_0_999 = 16'd-25509;
parameter WEIGHT_0_1000 = 16'd-2605;
parameter WEIGHT_0_1001 = 16'd1412;
parameter WEIGHT_0_1002 = 16'd4132;
parameter WEIGHT_0_1003 = 16'd6971;
parameter WEIGHT_0_1004 = 16'd-13494;
parameter WEIGHT_0_1005 = 16'd-29;
parameter WEIGHT_0_1006 = 16'd5163;
parameter WEIGHT_0_1007 = 16'd-14968;
parameter WEIGHT_0_1008 = 16'd-9480;
parameter WEIGHT_0_1009 = 16'd-23462;
parameter WEIGHT_0_1010 = 16'd-3853;
parameter WEIGHT_0_1011 = 16'd-8159;
parameter WEIGHT_0_1012 = 16'd2349;
parameter WEIGHT_0_1013 = 16'd6597;
parameter WEIGHT_0_1014 = 16'd-10707;
parameter WEIGHT_0_1015 = 16'd344;
parameter WEIGHT_0_1016 = 16'd5789;
parameter WEIGHT_0_1017 = 16'd-13333;
parameter WEIGHT_0_1018 = 16'd-10749;
parameter WEIGHT_0_1019 = 16'd-20096;
parameter WEIGHT_0_1020 = 16'd-13050;
parameter WEIGHT_0_1021 = 16'd-9587;
parameter WEIGHT_0_1022 = 16'd-3509;
parameter WEIGHT_0_1023 = 16'd5104;
parameter WEIGHT_0_1024 = 16'd-11164;
parameter WEIGHT_0_1025 = 16'd5982;
parameter WEIGHT_0_1026 = 16'd5903;
parameter WEIGHT_0_1027 = 16'd-8706;
parameter WEIGHT_0_1028 = 16'd-5232;
parameter WEIGHT_0_1029 = 16'd-13332;
parameter WEIGHT_0_1030 = 16'd-9188;
parameter WEIGHT_0_1031 = 16'd-9203;
parameter WEIGHT_0_1032 = 16'd-6192;
parameter WEIGHT_0_1033 = 16'd1983;
parameter WEIGHT_0_1034 = 16'd-5001;
parameter WEIGHT_0_1035 = 16'd2218;
parameter WEIGHT_0_1036 = 16'd5695;
parameter WEIGHT_0_1037 = 16'd-8184;
parameter WEIGHT_0_1038 = 16'd-11868;
parameter WEIGHT_0_1039 = 16'd-13688;
parameter WEIGHT_0_1040 = 16'd-7344;
parameter WEIGHT_0_1041 = 16'd-11480;
parameter WEIGHT_0_1042 = 16'd-6735;
parameter WEIGHT_0_1043 = 16'd1325;
parameter WEIGHT_0_1044 = 16'd-2536;
parameter WEIGHT_0_1045 = 16'd3635;
parameter WEIGHT_0_1046 = 16'd6481;
parameter WEIGHT_0_1047 = 16'd-6193;
parameter WEIGHT_0_1048 = 16'd-8746;
parameter WEIGHT_0_1049 = 16'd-16454;
parameter WEIGHT_0_1050 = 16'd-10788;
parameter WEIGHT_0_1051 = 16'd-6772;
parameter WEIGHT_0_1052 = 16'd-6478;
parameter WEIGHT_0_1053 = 16'd-3019;
parameter WEIGHT_0_1054 = 16'd-2114;
parameter WEIGHT_0_1055 = 16'd3420;
parameter WEIGHT_0_1056 = 16'd4105;
parameter WEIGHT_0_1057 = 16'd-5995;
parameter WEIGHT_0_1058 = 16'd-2769;
parameter WEIGHT_0_1059 = 16'd-13815;
parameter WEIGHT_0_1060 = 16'd-8134;
parameter WEIGHT_0_1061 = 16'd-12907;
parameter WEIGHT_0_1062 = 16'd-7931;
parameter WEIGHT_0_1063 = 16'd-11655;
parameter WEIGHT_0_1064 = 16'd-2231;
parameter WEIGHT_0_1065 = 16'd1520;
parameter WEIGHT_0_1066 = 16'd8948;
parameter WEIGHT_0_1067 = 16'd-5808;
parameter WEIGHT_0_1068 = 16'd-297;
parameter WEIGHT_0_1069 = 16'd-6464;
parameter WEIGHT_0_1070 = 16'd-7164;
parameter WEIGHT_0_1071 = 16'd-7991;
parameter WEIGHT_0_1072 = 16'd-15954;
parameter WEIGHT_0_1073 = 16'd-10595;
parameter WEIGHT_0_1074 = 16'd1118;
parameter WEIGHT_0_1075 = 16'd-361;
parameter WEIGHT_0_1076 = 16'd9214;
parameter WEIGHT_0_1077 = 16'd-64;
parameter WEIGHT_0_1078 = 16'd2075;
parameter WEIGHT_0_1079 = 16'd-869;
parameter WEIGHT_0_1080 = 16'd-3028;
parameter WEIGHT_0_1081 = 16'd-10417;
parameter WEIGHT_0_1082 = 16'd-4011;
parameter WEIGHT_0_1083 = 16'd-3328;
parameter WEIGHT_0_1084 = 16'd-7085;
parameter WEIGHT_0_1085 = 16'd481;
parameter WEIGHT_0_1086 = 16'd3221;
parameter WEIGHT_0_1087 = 16'd1435;
parameter WEIGHT_0_1088 = 16'd-445;
parameter WEIGHT_0_1089 = 16'd-5194;
parameter WEIGHT_0_1090 = 16'd-1693;
parameter WEIGHT_0_1091 = 16'd-3825;
parameter WEIGHT_0_1092 = 16'd1039;
parameter WEIGHT_0_1093 = 16'd-5208;
parameter WEIGHT_0_1094 = 16'd-5437;
parameter WEIGHT_0_1095 = 16'd-695;
parameter WEIGHT_0_1096 = 16'd2200;
parameter WEIGHT_0_1097 = 16'd-3046;
parameter WEIGHT_0_1098 = 16'd-2824;
parameter WEIGHT_0_1099 = 16'd-474;
parameter WEIGHT_0_1100 = 16'd-1940;
parameter WEIGHT_0_1101 = 16'd-5587;
parameter WEIGHT_0_1102 = 16'd-2726;
parameter WEIGHT_0_1103 = 16'd-444;
parameter WEIGHT_0_1104 = 16'd-274;
parameter WEIGHT_0_1105 = 16'd738;
parameter WEIGHT_0_1106 = 16'd2421;
parameter WEIGHT_0_1107 = 16'd-1468;
parameter WEIGHT_0_1108 = 16'd-5827;
parameter WEIGHT_0_1109 = 16'd-3362;
parameter WEIGHT_0_1110 = 16'd-1868;
parameter WEIGHT_0_1111 = 16'd-49;
parameter WEIGHT_0_1112 = 16'd-622;
parameter WEIGHT_0_1113 = 16'd-1958;
parameter WEIGHT_0_1114 = 16'd-501;
parameter WEIGHT_0_1115 = 16'd-529;
parameter WEIGHT_0_1116 = 16'd-853;
parameter WEIGHT_0_1117 = 16'd-388;
parameter WEIGHT_0_1118 = 16'd-1858;
parameter WEIGHT_0_1119 = 16'd1359;
parameter WEIGHT_0_1120 = 16'd332;
parameter WEIGHT_0_1121 = 16'd-501;
parameter WEIGHT_0_1122 = 16'd-1032;
parameter WEIGHT_0_1123 = 16'd2204;
parameter WEIGHT_0_1124 = 16'd1247;
parameter WEIGHT_0_1125 = 16'd2574;
parameter WEIGHT_0_1126 = 16'd2672;
parameter WEIGHT_0_1127 = 16'd-1848;
parameter WEIGHT_0_1128 = 16'd-1197;
parameter WEIGHT_0_1129 = 16'd575;
parameter WEIGHT_0_1130 = 16'd-485;
parameter WEIGHT_0_1131 = 16'd-1162;
parameter WEIGHT_0_1132 = 16'd-4807;
parameter WEIGHT_0_1133 = 16'd1320;
parameter WEIGHT_0_1134 = 16'd-762;
parameter WEIGHT_0_1135 = 16'd-725;
parameter WEIGHT_0_1136 = 16'd-1247;
parameter WEIGHT_0_1137 = 16'd1831;
parameter WEIGHT_0_1138 = 16'd-2821;
parameter WEIGHT_0_1139 = 16'd1257;
parameter WEIGHT_0_1140 = 16'd-3833;
parameter WEIGHT_0_1141 = 16'd-359;
parameter WEIGHT_0_1142 = 16'd-7245;
parameter WEIGHT_0_1143 = 16'd-1659;
parameter WEIGHT_0_1144 = 16'd-4592;
parameter WEIGHT_0_1145 = 16'd-4574;
parameter WEIGHT_0_1146 = 16'd-1230;
parameter WEIGHT_0_1147 = 16'd-1003;
parameter WEIGHT_0_1148 = 16'd223;
parameter WEIGHT_0_1149 = 16'd265;
parameter WEIGHT_0_1150 = 16'd1005;
parameter WEIGHT_0_1151 = 16'd-2631;
parameter WEIGHT_0_1152 = 16'd-2898;
parameter WEIGHT_0_1153 = 16'd3721;
parameter WEIGHT_0_1154 = 16'd-6776;
parameter WEIGHT_0_1155 = 16'd-3580;
parameter WEIGHT_0_1156 = 16'd-461;
parameter WEIGHT_0_1157 = 16'd484;
parameter WEIGHT_0_1158 = 16'd-8794;
parameter WEIGHT_0_1159 = 16'd-1993;
parameter WEIGHT_0_1160 = 16'd-8948;
parameter WEIGHT_0_1161 = 16'd1629;
parameter WEIGHT_0_1162 = 16'd-3029;
parameter WEIGHT_0_1163 = 16'd6649;
parameter WEIGHT_0_1164 = 16'd-517;
parameter WEIGHT_0_1165 = 16'd-11192;
parameter WEIGHT_0_1166 = 16'd3659;
parameter WEIGHT_0_1167 = 16'd-2705;
parameter WEIGHT_0_1168 = 16'd-9179;
parameter WEIGHT_0_1169 = 16'd-4912;
parameter WEIGHT_0_1170 = 16'd-7031;
parameter WEIGHT_0_1171 = 16'd-1777;
parameter WEIGHT_0_1172 = 16'd-1930;
parameter WEIGHT_0_1173 = 16'd7720;
parameter WEIGHT_0_1174 = 16'd2589;
parameter WEIGHT_0_1175 = 16'd-8844;
parameter WEIGHT_0_1176 = 16'd-1155;
parameter WEIGHT_0_1177 = 16'd-4863;
parameter WEIGHT_0_1178 = 16'd-11928;
parameter WEIGHT_0_1179 = 16'd-6622;
parameter WEIGHT_0_1180 = 16'd-5429;
parameter WEIGHT_0_1181 = 16'd-4149;
parameter WEIGHT_0_1182 = 16'd2397;
parameter WEIGHT_0_1183 = 16'd4384;
parameter WEIGHT_0_1184 = 16'd-4754;
parameter WEIGHT_0_1185 = 16'd-7655;
parameter WEIGHT_0_1186 = 16'd-195;
parameter WEIGHT_0_1187 = 16'd-7145;
parameter WEIGHT_0_1188 = 16'd-8587;
parameter WEIGHT_0_1189 = 16'd-5241;
parameter WEIGHT_0_1190 = 16'd-4472;
parameter WEIGHT_0_1191 = 16'd-3997;
parameter WEIGHT_0_1192 = 16'd806;
parameter WEIGHT_0_1193 = 16'd8481;
parameter WEIGHT_0_1194 = 16'd-2722;
parameter WEIGHT_0_1195 = 16'd-4287;
parameter WEIGHT_0_1196 = 16'd1531;
parameter WEIGHT_0_1197 = 16'd-10046;
parameter WEIGHT_0_1198 = 16'd-5640;
parameter WEIGHT_0_1199 = 16'd-7119;
parameter WEIGHT_0_1200 = 16'd-663;
parameter WEIGHT_0_1201 = 16'd-6796;
parameter WEIGHT_0_1202 = 16'd2858;
parameter WEIGHT_0_1203 = 16'd9178;
parameter WEIGHT_0_1204 = 16'd-8313;
parameter WEIGHT_0_1205 = 16'd-12999;
parameter WEIGHT_0_1206 = 16'd393;
parameter WEIGHT_0_1207 = 16'd-14469;
parameter WEIGHT_0_1208 = 16'd-2835;
parameter WEIGHT_0_1209 = 16'd-17467;
parameter WEIGHT_0_1210 = 16'd-3363;
parameter WEIGHT_0_1211 = 16'd-4634;
parameter WEIGHT_0_1212 = 16'd7465;
parameter WEIGHT_0_1213 = 16'd3514;
parameter WEIGHT_0_1214 = 16'd-9547;
parameter WEIGHT_0_1215 = 16'd-7561;
parameter WEIGHT_0_1216 = 16'd1851;
parameter WEIGHT_0_1217 = 16'd-17225;
parameter WEIGHT_0_1218 = 16'd904;
parameter WEIGHT_0_1219 = 16'd-20676;
parameter WEIGHT_0_1220 = 16'd-2538;
parameter WEIGHT_0_1221 = 16'd-2875;
parameter WEIGHT_0_1222 = 16'd7754;
parameter WEIGHT_0_1223 = 16'd8655;
parameter WEIGHT_0_1224 = 16'd-11505;
parameter WEIGHT_0_1225 = 16'd-3762;
parameter WEIGHT_0_1226 = 16'd1654;
parameter WEIGHT_0_1227 = 16'd-20114;
parameter WEIGHT_0_1228 = 16'd-2747;
parameter WEIGHT_0_1229 = 16'd-18021;
parameter WEIGHT_0_1230 = 16'd-801;
parameter WEIGHT_0_1231 = 16'd-6234;
parameter WEIGHT_0_1232 = 16'd4736;
parameter WEIGHT_0_1233 = 16'd6753;
parameter WEIGHT_0_1234 = 16'd-12928;
parameter WEIGHT_0_1235 = 16'd-1975;
parameter WEIGHT_0_1236 = 16'd-3084;
parameter WEIGHT_0_1237 = 16'd-14075;
parameter WEIGHT_0_1238 = 16'd-844;
parameter WEIGHT_0_1239 = 16'd-13908;
parameter WEIGHT_0_1240 = 16'd-1829;
parameter WEIGHT_0_1241 = 16'd543;
parameter WEIGHT_0_1242 = 16'd5178;
parameter WEIGHT_0_1243 = 16'd4969;
parameter WEIGHT_0_1244 = 16'd-9463;
parameter WEIGHT_0_1245 = 16'd-3348;
parameter WEIGHT_0_1246 = 16'd-6047;
parameter WEIGHT_0_1247 = 16'd-15052;
parameter WEIGHT_0_1248 = 16'd1996;
parameter WEIGHT_0_1249 = 16'd-13978;
parameter WEIGHT_0_1250 = 16'd-2287;
parameter WEIGHT_0_1251 = 16'd2228;
parameter WEIGHT_0_1252 = 16'd6831;
parameter WEIGHT_0_1253 = 16'd8212;
parameter WEIGHT_0_1254 = 16'd-6570;
parameter WEIGHT_0_1255 = 16'd-4430;
parameter WEIGHT_0_1256 = 16'd-612;
parameter WEIGHT_0_1257 = 16'd-16444;
parameter WEIGHT_0_1258 = 16'd899;
parameter WEIGHT_0_1259 = 16'd-8883;
parameter WEIGHT_0_1260 = 16'd107;
parameter WEIGHT_0_1261 = 16'd2325;
parameter WEIGHT_0_1262 = 16'd6720;
parameter WEIGHT_0_1263 = 16'd4956;
parameter WEIGHT_0_1264 = 16'd-10120;
parameter WEIGHT_0_1265 = 16'd-3164;
parameter WEIGHT_0_1266 = 16'd-3039;
parameter WEIGHT_0_1267 = 16'd-15233;
parameter WEIGHT_0_1268 = 16'd4677;
parameter WEIGHT_0_1269 = 16'd-13252;
parameter WEIGHT_0_1270 = 16'd-5;
parameter WEIGHT_0_1271 = 16'd1644;
parameter WEIGHT_0_1272 = 16'd1929;
parameter WEIGHT_0_1273 = 16'd6680;
parameter WEIGHT_0_1274 = 16'd-12629;
parameter WEIGHT_0_1275 = 16'd2284;
parameter WEIGHT_0_1276 = 16'd-3342;
parameter WEIGHT_0_1277 = 16'd-15231;
parameter WEIGHT_0_1278 = 16'd3713;
parameter WEIGHT_0_1279 = 16'd-16132;
parameter WEIGHT_0_1280 = 16'd-2181;
parameter WEIGHT_0_1281 = 16'd412;
parameter WEIGHT_0_1282 = 16'd3184;
parameter WEIGHT_0_1283 = 16'd4187;
parameter WEIGHT_0_1284 = 16'd-4609;
parameter WEIGHT_0_1285 = 16'd2125;
parameter WEIGHT_0_1286 = 16'd-551;
parameter WEIGHT_0_1287 = 16'd-17192;
parameter WEIGHT_0_1288 = 16'd2635;
parameter WEIGHT_0_1289 = 16'd-18501;
parameter WEIGHT_0_1290 = 16'd995;
parameter WEIGHT_0_1291 = 16'd-659;
parameter WEIGHT_0_1292 = 16'd514;
parameter WEIGHT_0_1293 = 16'd1928;
parameter WEIGHT_0_1294 = 16'd-3766;
parameter WEIGHT_0_1295 = 16'd5812;
parameter WEIGHT_0_1296 = 16'd3844;
parameter WEIGHT_0_1297 = 16'd-20718;
parameter WEIGHT_0_1298 = 16'd48;
parameter WEIGHT_0_1299 = 16'd-17030;
parameter WEIGHT_0_1300 = 16'd-2652;
parameter WEIGHT_0_1301 = 16'd-541;
parameter WEIGHT_0_1302 = 16'd-1835;
parameter WEIGHT_0_1303 = 16'd2501;
parameter WEIGHT_0_1304 = 16'd-4167;
parameter WEIGHT_0_1305 = 16'd3447;
parameter WEIGHT_0_1306 = 16'd3858;
parameter WEIGHT_0_1307 = 16'd-18146;
parameter WEIGHT_0_1308 = 16'd-82;
parameter WEIGHT_0_1309 = 16'd-15930;
parameter WEIGHT_0_1310 = 16'd-4601;
parameter WEIGHT_0_1311 = 16'd3001;
parameter WEIGHT_0_1312 = 16'd-3265;
parameter WEIGHT_0_1313 = 16'd1296;
parameter WEIGHT_0_1314 = 16'd412;
parameter WEIGHT_0_1315 = 16'd1522;
parameter WEIGHT_0_1316 = 16'd6176;
parameter WEIGHT_0_1317 = 16'd-13537;
parameter WEIGHT_0_1318 = 16'd-2713;
parameter WEIGHT_0_1319 = 16'd-15067;
parameter WEIGHT_0_1320 = 16'd-1944;
parameter WEIGHT_0_1321 = 16'd1514;
parameter WEIGHT_0_1322 = 16'd-4043;
parameter WEIGHT_0_1323 = 16'd-5756;
parameter WEIGHT_0_1324 = 16'd3568;
parameter WEIGHT_0_1325 = 16'd-591;
parameter WEIGHT_0_1326 = 16'd7437;
parameter WEIGHT_0_1327 = 16'd-13520;
parameter WEIGHT_0_1328 = 16'd-346;
parameter WEIGHT_0_1329 = 16'd-15339;
parameter WEIGHT_0_1330 = 16'd-2857;
parameter WEIGHT_0_1331 = 16'd1784;
parameter WEIGHT_0_1332 = 16'd-10289;
parameter WEIGHT_0_1333 = 16'd-6546;
parameter WEIGHT_0_1334 = 16'd3995;
parameter WEIGHT_0_1335 = 16'd1718;
parameter WEIGHT_0_1336 = 16'd8382;
parameter WEIGHT_0_1337 = 16'd-7917;
parameter WEIGHT_0_1338 = 16'd-3321;
parameter WEIGHT_0_1339 = 16'd-25029;
parameter WEIGHT_0_1340 = 16'd-4925;
parameter WEIGHT_0_1341 = 16'd-1643;
parameter WEIGHT_0_1342 = 16'd-11102;
parameter WEIGHT_0_1343 = 16'd-10587;
parameter WEIGHT_0_1344 = 16'd3448;
parameter WEIGHT_0_1345 = 16'd1336;
parameter WEIGHT_0_1346 = 16'd11538;
parameter WEIGHT_0_1347 = 16'd-9467;
parameter WEIGHT_0_1348 = 16'd-4250;
parameter WEIGHT_0_1349 = 16'd-16263;
parameter WEIGHT_0_1350 = 16'd-3655;
parameter WEIGHT_0_1351 = 16'd483;
parameter WEIGHT_0_1352 = 16'd-15764;
parameter WEIGHT_0_1353 = 16'd-17857;
parameter WEIGHT_0_1354 = 16'd4401;
parameter WEIGHT_0_1355 = 16'd3005;
parameter WEIGHT_0_1356 = 16'd5883;
parameter WEIGHT_0_1357 = 16'd-6598;
parameter WEIGHT_0_1358 = 16'd-5563;
parameter WEIGHT_0_1359 = 16'd-12039;
parameter WEIGHT_0_1360 = 16'd-8493;
parameter WEIGHT_0_1361 = 16'd-10462;
parameter WEIGHT_0_1362 = 16'd-11251;
parameter WEIGHT_0_1363 = 16'd-16981;
parameter WEIGHT_0_1364 = 16'd2591;
parameter WEIGHT_0_1365 = 16'd7372;
parameter WEIGHT_0_1366 = 16'd3163;
parameter WEIGHT_0_1367 = 16'd-7559;
parameter WEIGHT_0_1368 = 16'd-2120;
parameter WEIGHT_0_1369 = 16'd-8514;
parameter WEIGHT_0_1370 = 16'd-9941;
parameter WEIGHT_0_1371 = 16'd-14112;
parameter WEIGHT_0_1372 = 16'd140;
parameter WEIGHT_0_1373 = 16'd-5037;
parameter WEIGHT_0_1374 = 16'd-975;
parameter WEIGHT_0_1375 = 16'd7987;
parameter WEIGHT_0_1376 = 16'd2358;
parameter WEIGHT_0_1377 = 16'd-5586;
parameter WEIGHT_0_1378 = 16'd2762;
parameter WEIGHT_0_1379 = 16'd-5305;
parameter WEIGHT_0_1380 = 16'd-7584;
parameter WEIGHT_0_1381 = 16'd-4703;
parameter WEIGHT_0_1382 = 16'd-3711;
parameter WEIGHT_0_1383 = 16'd-1316;
parameter WEIGHT_0_1384 = 16'd-4902;
parameter WEIGHT_0_1385 = 16'd2005;
parameter WEIGHT_0_1386 = 16'd-1672;
parameter WEIGHT_0_1387 = 16'd-2642;
parameter WEIGHT_0_1388 = 16'd634;
parameter WEIGHT_0_1389 = 16'd-3550;
parameter WEIGHT_0_1390 = 16'd154;
parameter WEIGHT_0_1391 = 16'd-4174;
parameter WEIGHT_0_1392 = 16'd-4238;
parameter WEIGHT_0_1393 = 16'd930;
parameter WEIGHT_0_1394 = 16'd-3979;
parameter WEIGHT_0_1395 = 16'd-4912;
parameter WEIGHT_0_1396 = 16'd404;
parameter WEIGHT_0_1397 = 16'd-1293;
parameter WEIGHT_0_1398 = 16'd1384;
parameter WEIGHT_0_1399 = 16'd-3409;
parameter WEIGHT_0_1400 = 16'd-126;
parameter WEIGHT_0_1401 = 16'd-2583;
parameter WEIGHT_0_1402 = 16'd613;
parameter WEIGHT_0_1403 = 16'd-367;
parameter WEIGHT_0_1404 = 16'd-1060;
parameter WEIGHT_0_1405 = 16'd-384;
parameter WEIGHT_0_1406 = 16'd1167;
parameter WEIGHT_0_1407 = 16'd687;
parameter WEIGHT_0_1408 = 16'd-2661;
parameter WEIGHT_0_1409 = 16'd-545;
parameter WEIGHT_0_1410 = 16'd1670;
parameter WEIGHT_0_1411 = 16'd-1279;
parameter WEIGHT_0_1412 = 16'd-219;
parameter WEIGHT_0_1413 = 16'd-2535;
parameter WEIGHT_0_1414 = 16'd-743;
parameter WEIGHT_0_1415 = 16'd1797;
parameter WEIGHT_0_1416 = 16'd92;
parameter WEIGHT_0_1417 = 16'd2012;
parameter WEIGHT_0_1418 = 16'd-737;
parameter WEIGHT_0_1419 = 16'd-2726;
parameter WEIGHT_0_1420 = 16'd-5026;
parameter WEIGHT_0_1421 = 16'd607;
parameter WEIGHT_0_1422 = 16'd2806;
parameter WEIGHT_0_1423 = 16'd-372;
parameter WEIGHT_0_1424 = 16'd-2574;
parameter WEIGHT_0_1425 = 16'd-2723;
parameter WEIGHT_0_1426 = 16'd1508;
parameter WEIGHT_0_1427 = 16'd-3418;
parameter WEIGHT_0_1428 = 16'd-3332;
parameter WEIGHT_0_1429 = 16'd-5472;
parameter WEIGHT_0_1430 = 16'd-1414;
parameter WEIGHT_0_1431 = 16'd3133;
parameter WEIGHT_0_1432 = 16'd-2978;
parameter WEIGHT_0_1433 = 16'd4318;
parameter WEIGHT_0_1434 = 16'd-658;
parameter WEIGHT_0_1435 = 16'd-7263;
parameter WEIGHT_0_1436 = 16'd-4340;
parameter WEIGHT_0_1437 = 16'd-1545;
parameter WEIGHT_0_1438 = 16'd-5345;
parameter WEIGHT_0_1439 = 16'd-5322;
parameter WEIGHT_0_1440 = 16'd-10124;
parameter WEIGHT_0_1441 = 16'd1728;
parameter WEIGHT_0_1442 = 16'd1717;
parameter WEIGHT_0_1443 = 16'd9756;
parameter WEIGHT_0_1444 = 16'd3145;
parameter WEIGHT_0_1445 = 16'd-12966;
parameter WEIGHT_0_1446 = 16'd-1819;
parameter WEIGHT_0_1447 = 16'd-5969;
parameter WEIGHT_0_1448 = 16'd-9824;
parameter WEIGHT_0_1449 = 16'd-2982;
parameter WEIGHT_0_1450 = 16'd-8819;
parameter WEIGHT_0_1451 = 16'd1920;
parameter WEIGHT_0_1452 = 16'd2387;
parameter WEIGHT_0_1453 = 16'd9252;
parameter WEIGHT_0_1454 = 16'd3451;
parameter WEIGHT_0_1455 = 16'd-11386;
parameter WEIGHT_0_1456 = 16'd-4102;
parameter WEIGHT_0_1457 = 16'd-919;
parameter WEIGHT_0_1458 = 16'd-11477;
parameter WEIGHT_0_1459 = 16'd-10757;
parameter WEIGHT_0_1460 = 16'd-6740;
parameter WEIGHT_0_1461 = 16'd-2901;
parameter WEIGHT_0_1462 = 16'd3369;
parameter WEIGHT_0_1463 = 16'd9534;
parameter WEIGHT_0_1464 = 16'd3187;
parameter WEIGHT_0_1465 = 16'd-9516;
parameter WEIGHT_0_1466 = 16'd-1318;
parameter WEIGHT_0_1467 = 16'd683;
parameter WEIGHT_0_1468 = 16'd-9306;
parameter WEIGHT_0_1469 = 16'd-20632;
parameter WEIGHT_0_1470 = 16'd-1848;
parameter WEIGHT_0_1471 = 16'd-6617;
parameter WEIGHT_0_1472 = 16'd2781;
parameter WEIGHT_0_1473 = 16'd3428;
parameter WEIGHT_0_1474 = 16'd-2475;
parameter WEIGHT_0_1475 = 16'd-6175;
parameter WEIGHT_0_1476 = 16'd-3389;
parameter WEIGHT_0_1477 = 16'd296;
parameter WEIGHT_0_1478 = 16'd-5000;
parameter WEIGHT_0_1479 = 16'd-16463;
parameter WEIGHT_0_1480 = 16'd-3116;
parameter WEIGHT_0_1481 = 16'd-9496;
parameter WEIGHT_0_1482 = 16'd5422;
parameter WEIGHT_0_1483 = 16'd3118;
parameter WEIGHT_0_1484 = 16'd-1911;
parameter WEIGHT_0_1485 = 16'd-1546;
parameter WEIGHT_0_1486 = 16'd1267;
parameter WEIGHT_0_1487 = 16'd556;
parameter WEIGHT_0_1488 = 16'd-3063;
parameter WEIGHT_0_1489 = 16'd-10787;
parameter WEIGHT_0_1490 = 16'd-2138;
parameter WEIGHT_0_1491 = 16'd-7916;
parameter WEIGHT_0_1492 = 16'd4387;
parameter WEIGHT_0_1493 = 16'd6265;
parameter WEIGHT_0_1494 = 16'd-1976;
parameter WEIGHT_0_1495 = 16'd-1039;
parameter WEIGHT_0_1496 = 16'd-1579;
parameter WEIGHT_0_1497 = 16'd-821;
parameter WEIGHT_0_1498 = 16'd-3568;
parameter WEIGHT_0_1499 = 16'd-12548;
parameter WEIGHT_0_1500 = 16'd-1141;
parameter WEIGHT_0_1501 = 16'd-6998;
parameter WEIGHT_0_1502 = 16'd4134;
parameter WEIGHT_0_1503 = 16'd3290;
parameter WEIGHT_0_1504 = 16'd-5607;
parameter WEIGHT_0_1505 = 16'd1423;
parameter WEIGHT_0_1506 = 16'd-1203;
parameter WEIGHT_0_1507 = 16'd-3546;
parameter WEIGHT_0_1508 = 16'd-3472;
parameter WEIGHT_0_1509 = 16'd-3731;
parameter WEIGHT_0_1510 = 16'd-2853;
parameter WEIGHT_0_1511 = 16'd-3954;
parameter WEIGHT_0_1512 = 16'd7876;
parameter WEIGHT_0_1513 = 16'd4513;
parameter WEIGHT_0_1514 = 16'd-3439;
parameter WEIGHT_0_1515 = 16'd-2299;
parameter WEIGHT_0_1516 = 16'd-5646;
parameter WEIGHT_0_1517 = 16'd-6690;
parameter WEIGHT_0_1518 = 16'd-220;
parameter WEIGHT_0_1519 = 16'd755;
parameter WEIGHT_0_1520 = 16'd-2676;
parameter WEIGHT_0_1521 = 16'd-1812;
parameter WEIGHT_0_1522 = 16'd3649;
parameter WEIGHT_0_1523 = 16'd1503;
parameter WEIGHT_0_1524 = 16'd-4798;
parameter WEIGHT_0_1525 = 16'd-1917;
parameter WEIGHT_0_1526 = 16'd-4532;
parameter WEIGHT_0_1527 = 16'd-7941;
parameter WEIGHT_0_1528 = 16'd5281;
parameter WEIGHT_0_1529 = 16'd531;
parameter WEIGHT_0_1530 = 16'd2668;
parameter WEIGHT_0_1531 = 16'd-1894;
parameter WEIGHT_0_1532 = 16'd4734;
parameter WEIGHT_0_1533 = 16'd3077;
parameter WEIGHT_0_1534 = 16'd-8319;
parameter WEIGHT_0_1535 = 16'd-230;
parameter WEIGHT_0_1536 = 16'd-4939;
parameter WEIGHT_0_1537 = 16'd-10222;
parameter WEIGHT_0_1538 = 16'd2779;
parameter WEIGHT_0_1539 = 16'd-2107;
parameter WEIGHT_0_1540 = 16'd1070;
parameter WEIGHT_0_1541 = 16'd-124;
parameter WEIGHT_0_1542 = 16'd3503;
parameter WEIGHT_0_1543 = 16'd1212;
parameter WEIGHT_0_1544 = 16'd-1667;
parameter WEIGHT_0_1545 = 16'd-5386;
parameter WEIGHT_0_1546 = 16'd-5164;
parameter WEIGHT_0_1547 = 16'd-9694;
parameter WEIGHT_0_1548 = 16'd3933;
parameter WEIGHT_0_1549 = 16'd-6836;
parameter WEIGHT_0_1550 = 16'd4436;
parameter WEIGHT_0_1551 = 16'd-671;
parameter WEIGHT_0_1552 = 16'd6637;
parameter WEIGHT_0_1553 = 16'd2248;
parameter WEIGHT_0_1554 = 16'd-2245;
parameter WEIGHT_0_1555 = 16'd-1402;
parameter WEIGHT_0_1556 = 16'd-713;
parameter WEIGHT_0_1557 = 16'd-12592;
parameter WEIGHT_0_1558 = 16'd5355;
parameter WEIGHT_0_1559 = 16'd-8056;
parameter WEIGHT_0_1560 = 16'd3788;
parameter WEIGHT_0_1561 = 16'd-4317;
parameter WEIGHT_0_1562 = 16'd7297;
parameter WEIGHT_0_1563 = 16'd2428;
parameter WEIGHT_0_1564 = 16'd445;
parameter WEIGHT_0_1565 = 16'd30;
parameter WEIGHT_0_1566 = 16'd-3798;
parameter WEIGHT_0_1567 = 16'd-11107;
parameter WEIGHT_0_1568 = 16'd4832;
parameter WEIGHT_0_1569 = 16'd-10276;
parameter WEIGHT_0_1570 = 16'd3925;
parameter WEIGHT_0_1571 = 16'd-6396;
parameter WEIGHT_0_1572 = 16'd6357;
parameter WEIGHT_0_1573 = 16'd-1194;
parameter WEIGHT_0_1574 = 16'd-1667;
parameter WEIGHT_0_1575 = 16'd1926;
parameter WEIGHT_0_1576 = 16'd-300;
parameter WEIGHT_0_1577 = 16'd-13097;
parameter WEIGHT_0_1578 = 16'd3399;
parameter WEIGHT_0_1579 = 16'd-13483;
parameter WEIGHT_0_1580 = 16'd4093;
parameter WEIGHT_0_1581 = 16'd-2588;
parameter WEIGHT_0_1582 = 16'd3276;
parameter WEIGHT_0_1583 = 16'd639;
parameter WEIGHT_0_1584 = 16'd2212;
parameter WEIGHT_0_1585 = 16'd1540;
parameter WEIGHT_0_1586 = 16'd828;
parameter WEIGHT_0_1587 = 16'd-16531;
parameter WEIGHT_0_1588 = 16'd-832;
parameter WEIGHT_0_1589 = 16'd-13060;
parameter WEIGHT_0_1590 = 16'd735;
parameter WEIGHT_0_1591 = 16'd709;
parameter WEIGHT_0_1592 = 16'd-900;
parameter WEIGHT_0_1593 = 16'd-3285;
parameter WEIGHT_0_1594 = 16'd2681;
parameter WEIGHT_0_1595 = 16'd2825;
parameter WEIGHT_0_1596 = 16'd4565;
parameter WEIGHT_0_1597 = 16'd-15809;
parameter WEIGHT_0_1598 = 16'd2316;
parameter WEIGHT_0_1599 = 16'd-8876;
parameter WEIGHT_0_1600 = 16'd750;
parameter WEIGHT_0_1601 = 16'd3508;
parameter WEIGHT_0_1602 = 16'd-1970;
parameter WEIGHT_0_1603 = 16'd-2925;
parameter WEIGHT_0_1604 = 16'd1351;
parameter WEIGHT_0_1605 = 16'd3090;
parameter WEIGHT_0_1606 = 16'd5139;
parameter WEIGHT_0_1607 = 16'd-21333;
parameter WEIGHT_0_1608 = 16'd3061;
parameter WEIGHT_0_1609 = 16'd-10362;
parameter WEIGHT_0_1610 = 16'd-1042;
parameter WEIGHT_0_1611 = 16'd6195;
parameter WEIGHT_0_1612 = 16'd31;
parameter WEIGHT_0_1613 = 16'd-6393;
parameter WEIGHT_0_1614 = 16'd3497;
parameter WEIGHT_0_1615 = 16'd3446;
parameter WEIGHT_0_1616 = 16'd6027;
parameter WEIGHT_0_1617 = 16'd-15770;
parameter WEIGHT_0_1618 = 16'd622;
parameter WEIGHT_0_1619 = 16'd-14903;
parameter WEIGHT_0_1620 = 16'd-1826;
parameter WEIGHT_0_1621 = 16'd4075;
parameter WEIGHT_0_1622 = 16'd-3822;
parameter WEIGHT_0_1623 = 16'd-8622;
parameter WEIGHT_0_1624 = 16'd6860;
parameter WEIGHT_0_1625 = 16'd5781;
parameter WEIGHT_0_1626 = 16'd6539;
parameter WEIGHT_0_1627 = 16'd-13631;
parameter WEIGHT_0_1628 = 16'd-3863;
parameter WEIGHT_0_1629 = 16'd-16789;
parameter WEIGHT_0_1630 = 16'd-6425;
parameter WEIGHT_0_1631 = 16'd4039;
parameter WEIGHT_0_1632 = 16'd-11512;
parameter WEIGHT_0_1633 = 16'd-12021;
parameter WEIGHT_0_1634 = 16'd10338;
parameter WEIGHT_0_1635 = 16'd5093;
parameter WEIGHT_0_1636 = 16'd6751;
parameter WEIGHT_0_1637 = 16'd-18647;
parameter WEIGHT_0_1638 = 16'd-7564;
parameter WEIGHT_0_1639 = 16'd-24523;
parameter WEIGHT_0_1640 = 16'd-8103;
parameter WEIGHT_0_1641 = 16'd-2796;
parameter WEIGHT_0_1642 = 16'd-15841;
parameter WEIGHT_0_1643 = 16'd-14077;
parameter WEIGHT_0_1644 = 16'd4009;
parameter WEIGHT_0_1645 = 16'd8025;
parameter WEIGHT_0_1646 = 16'd4525;
parameter WEIGHT_0_1647 = 16'd-13151;
parameter WEIGHT_0_1648 = 16'd-5076;
parameter WEIGHT_0_1649 = 16'd-18983;
parameter WEIGHT_0_1650 = 16'd-17181;
parameter WEIGHT_0_1651 = 16'd-12284;
parameter WEIGHT_0_1652 = 16'd-5498;
parameter WEIGHT_0_1653 = 16'd-14739;
parameter WEIGHT_0_1654 = 16'd-1606;
parameter WEIGHT_0_1655 = 16'd8760;
parameter WEIGHT_0_1656 = 16'd1222;
parameter WEIGHT_0_1657 = 16'd-6551;
parameter WEIGHT_0_1658 = 16'd1413;
parameter WEIGHT_0_1659 = 16'd-14034;
parameter WEIGHT_0_1660 = 16'd-14716;
parameter WEIGHT_0_1661 = 16'd-8291;
parameter WEIGHT_0_1662 = 16'd-8085;
parameter WEIGHT_0_1663 = 16'd-9615;
parameter WEIGHT_0_1664 = 16'd-6446;
parameter WEIGHT_0_1665 = 16'd10006;
parameter WEIGHT_0_1666 = 16'd1083;
parameter WEIGHT_0_1667 = 16'd-5127;
parameter WEIGHT_0_1668 = 16'd-59;
parameter WEIGHT_0_1669 = 16'd-5327;
parameter WEIGHT_0_1670 = 16'd-4261;
parameter WEIGHT_0_1671 = 16'd-3016;
parameter WEIGHT_0_1672 = 16'd-2470;
parameter WEIGHT_0_1673 = 16'd-4849;
parameter WEIGHT_0_1674 = 16'd-3755;
parameter WEIGHT_0_1675 = 16'd1576;
parameter WEIGHT_0_1676 = 16'd280;
parameter WEIGHT_0_1677 = 16'd-2821;
parameter WEIGHT_0_1678 = 16'd-3067;
parameter WEIGHT_0_1679 = 16'd1241;
parameter WEIGHT_0_1680 = 16'd2525;
parameter WEIGHT_0_1681 = 16'd-549;
parameter WEIGHT_0_1682 = 16'd593;
parameter WEIGHT_0_1683 = 16'd600;
parameter WEIGHT_0_1684 = 16'd-185;
parameter WEIGHT_0_1685 = 16'd118;
parameter WEIGHT_0_1686 = 16'd-1948;
parameter WEIGHT_0_1687 = 16'd-1684;
parameter WEIGHT_0_1688 = 16'd55;
parameter WEIGHT_0_1689 = 16'd-2141;
parameter WEIGHT_0_1690 = 16'd-2404;
parameter WEIGHT_0_1691 = 16'd-2183;
parameter WEIGHT_0_1692 = 16'd-593;
parameter WEIGHT_0_1693 = 16'd5186;
parameter WEIGHT_0_1694 = 16'd-1317;
parameter WEIGHT_0_1695 = 16'd-3810;
parameter WEIGHT_0_1696 = 16'd-679;
parameter WEIGHT_0_1697 = 16'd-1167;
parameter WEIGHT_0_1698 = 16'd-4679;
parameter WEIGHT_0_1699 = 16'd-1393;
parameter WEIGHT_0_1700 = 16'd-4352;
parameter WEIGHT_0_1701 = 16'd-4848;
parameter WEIGHT_0_1702 = 16'd930;
parameter WEIGHT_0_1703 = 16'd507;
parameter WEIGHT_0_1704 = 16'd-2024;
parameter WEIGHT_0_1705 = 16'd-1286;
parameter WEIGHT_0_1706 = 16'd-1722;
parameter WEIGHT_0_1707 = 16'd4182;
parameter WEIGHT_0_1708 = 16'd-7163;
parameter WEIGHT_0_1709 = 16'd-6566;
parameter WEIGHT_0_1710 = 16'd-7609;
parameter WEIGHT_0_1711 = 16'd1737;
parameter WEIGHT_0_1712 = 16'd-3330;
parameter WEIGHT_0_1713 = 16'd6905;
parameter WEIGHT_0_1714 = 16'd-3583;
parameter WEIGHT_0_1715 = 16'd-8951;
parameter WEIGHT_0_1716 = 16'd-7445;
parameter WEIGHT_0_1717 = 16'd7171;
parameter WEIGHT_0_1718 = 16'd-6502;
parameter WEIGHT_0_1719 = 16'd-6109;
parameter WEIGHT_0_1720 = 16'd-11387;
parameter WEIGHT_0_1721 = 16'd2097;
parameter WEIGHT_0_1722 = 16'd2129;
parameter WEIGHT_0_1723 = 16'd7281;
parameter WEIGHT_0_1724 = 16'd1803;
parameter WEIGHT_0_1725 = 16'd-10063;
parameter WEIGHT_0_1726 = 16'd-3631;
parameter WEIGHT_0_1727 = 16'd1433;
parameter WEIGHT_0_1728 = 16'd-8856;
parameter WEIGHT_0_1729 = 16'd-11069;
parameter WEIGHT_0_1730 = 16'd-3071;
parameter WEIGHT_0_1731 = 16'd-5061;
parameter WEIGHT_0_1732 = 16'd3545;
parameter WEIGHT_0_1733 = 16'd3953;
parameter WEIGHT_0_1734 = 16'd5403;
parameter WEIGHT_0_1735 = 16'd-7675;
parameter WEIGHT_0_1736 = 16'd-5330;
parameter WEIGHT_0_1737 = 16'd2291;
parameter WEIGHT_0_1738 = 16'd-4741;
parameter WEIGHT_0_1739 = 16'd-17262;
parameter WEIGHT_0_1740 = 16'd-1472;
parameter WEIGHT_0_1741 = 16'd-1535;
parameter WEIGHT_0_1742 = 16'd3907;
parameter WEIGHT_0_1743 = 16'd5008;
parameter WEIGHT_0_1744 = 16'd-257;
parameter WEIGHT_0_1745 = 16'd-6006;
parameter WEIGHT_0_1746 = 16'd-8300;
parameter WEIGHT_0_1747 = 16'd4999;
parameter WEIGHT_0_1748 = 16'd-6264;
parameter WEIGHT_0_1749 = 16'd-15716;
parameter WEIGHT_0_1750 = 16'd-570;
parameter WEIGHT_0_1751 = 16'd-7757;
parameter WEIGHT_0_1752 = 16'd1840;
parameter WEIGHT_0_1753 = 16'd1342;
parameter WEIGHT_0_1754 = 16'd832;
parameter WEIGHT_0_1755 = 16'd-2755;
parameter WEIGHT_0_1756 = 16'd378;
parameter WEIGHT_0_1757 = 16'd4451;
parameter WEIGHT_0_1758 = 16'd-3023;
parameter WEIGHT_0_1759 = 16'd-14264;
parameter WEIGHT_0_1760 = 16'd-5870;
parameter WEIGHT_0_1761 = 16'd-8325;
parameter WEIGHT_0_1762 = 16'd3604;
parameter WEIGHT_0_1763 = 16'd3245;
parameter WEIGHT_0_1764 = 16'd1322;
parameter WEIGHT_0_1765 = 16'd-601;
parameter WEIGHT_0_1766 = 16'd-3505;
parameter WEIGHT_0_1767 = 16'd3593;
parameter WEIGHT_0_1768 = 16'd67;
parameter WEIGHT_0_1769 = 16'd-7980;
parameter WEIGHT_0_1770 = 16'd-4605;
parameter WEIGHT_0_1771 = 16'd-12947;
parameter WEIGHT_0_1772 = 16'd4447;
parameter WEIGHT_0_1773 = 16'd4364;
parameter WEIGHT_0_1774 = 16'd-2063;
parameter WEIGHT_0_1775 = 16'd-1645;
parameter WEIGHT_0_1776 = 16'd-645;
parameter WEIGHT_0_1777 = 16'd4053;
parameter WEIGHT_0_1778 = 16'd-2944;
parameter WEIGHT_0_1779 = 16'd-5300;
parameter WEIGHT_0_1780 = 16'd-576;
parameter WEIGHT_0_1781 = 16'd-8633;
parameter WEIGHT_0_1782 = 16'd542;
parameter WEIGHT_0_1783 = 16'd3109;
parameter WEIGHT_0_1784 = 16'd-4789;
parameter WEIGHT_0_1785 = 16'd1670;
parameter WEIGHT_0_1786 = 16'd-7029;
parameter WEIGHT_0_1787 = 16'd2462;
parameter WEIGHT_0_1788 = 16'd-912;
parameter WEIGHT_0_1789 = 16'd-1409;
parameter WEIGHT_0_1790 = 16'd-247;
parameter WEIGHT_0_1791 = 16'd-5142;
parameter WEIGHT_0_1792 = 16'd-731;
parameter WEIGHT_0_1793 = 16'd3396;
parameter WEIGHT_0_1794 = 16'd-5930;
parameter WEIGHT_0_1795 = 16'd1154;
parameter WEIGHT_0_1796 = 16'd-8624;
parameter WEIGHT_0_1797 = 16'd5594;
parameter WEIGHT_0_1798 = 16'd-2603;
parameter WEIGHT_0_1799 = 16'd-280;
parameter WEIGHT_0_1800 = 16'd135;
parameter WEIGHT_0_1801 = 16'd-5470;
parameter WEIGHT_0_1802 = 16'd2454;
parameter WEIGHT_0_1803 = 16'd2930;
parameter WEIGHT_0_1804 = 16'd-9104;
parameter WEIGHT_0_1805 = 16'd735;
parameter WEIGHT_0_1806 = 16'd-3182;
parameter WEIGHT_0_1807 = 16'd-1309;
parameter WEIGHT_0_1808 = 16'd3805;
parameter WEIGHT_0_1809 = 16'd4759;
parameter WEIGHT_0_1810 = 16'd4035;
parameter WEIGHT_0_1811 = 16'd-4122;
parameter WEIGHT_0_1812 = 16'd3870;
parameter WEIGHT_0_1813 = 16'd2186;
parameter WEIGHT_0_1814 = 16'd-11151;
parameter WEIGHT_0_1815 = 16'd991;
parameter WEIGHT_0_1816 = 16'd-6007;
parameter WEIGHT_0_1817 = 16'd-5100;
parameter WEIGHT_0_1818 = 16'd-896;
parameter WEIGHT_0_1819 = 16'd5248;
parameter WEIGHT_0_1820 = 16'd1798;
parameter WEIGHT_0_1821 = 16'd-7471;
parameter WEIGHT_0_1822 = 16'd880;
parameter WEIGHT_0_1823 = 16'd3929;
parameter WEIGHT_0_1824 = 16'd-10096;
parameter WEIGHT_0_1825 = 16'd2218;
parameter WEIGHT_0_1826 = 16'd-5157;
parameter WEIGHT_0_1827 = 16'd-2747;
parameter WEIGHT_0_1828 = 16'd3698;
parameter WEIGHT_0_1829 = 16'd9254;
parameter WEIGHT_0_1830 = 16'd4038;
parameter WEIGHT_0_1831 = 16'd-6753;
parameter WEIGHT_0_1832 = 16'd4110;
parameter WEIGHT_0_1833 = 16'd5864;
parameter WEIGHT_0_1834 = 16'd-12802;
parameter WEIGHT_0_1835 = 16'd-2768;
parameter WEIGHT_0_1836 = 16'd-3152;
parameter WEIGHT_0_1837 = 16'd-3358;
parameter WEIGHT_0_1838 = 16'd2276;
parameter WEIGHT_0_1839 = 16'd5116;
parameter WEIGHT_0_1840 = 16'd5970;
parameter WEIGHT_0_1841 = 16'd-6997;
parameter WEIGHT_0_1842 = 16'd4052;
parameter WEIGHT_0_1843 = 16'd4690;
parameter WEIGHT_0_1844 = 16'd-10512;
parameter WEIGHT_0_1845 = 16'd508;
parameter WEIGHT_0_1846 = 16'd-3045;
parameter WEIGHT_0_1847 = 16'd-569;
parameter WEIGHT_0_1848 = 16'd4396;
parameter WEIGHT_0_1849 = 16'd8009;
parameter WEIGHT_0_1850 = 16'd3798;
parameter WEIGHT_0_1851 = 16'd-7711;
parameter WEIGHT_0_1852 = 16'd-809;
parameter WEIGHT_0_1853 = 16'd2170;
parameter WEIGHT_0_1854 = 16'd-6670;
parameter WEIGHT_0_1855 = 16'd1151;
parameter WEIGHT_0_1856 = 16'd-1601;
parameter WEIGHT_0_1857 = 16'd-3967;
parameter WEIGHT_0_1858 = 16'd2546;
parameter WEIGHT_0_1859 = 16'd5601;
parameter WEIGHT_0_1860 = 16'd4276;
parameter WEIGHT_0_1861 = 16'd-3254;
parameter WEIGHT_0_1862 = 16'd689;
parameter WEIGHT_0_1863 = 16'd2426;
parameter WEIGHT_0_1864 = 16'd-6266;
parameter WEIGHT_0_1865 = 16'd2836;
parameter WEIGHT_0_1866 = 16'd-2073;
parameter WEIGHT_0_1867 = 16'd-3137;
parameter WEIGHT_0_1868 = 16'd2371;
parameter WEIGHT_0_1869 = 16'd3437;
parameter WEIGHT_0_1870 = 16'd2035;
parameter WEIGHT_0_1871 = 16'd-187;
parameter WEIGHT_0_1872 = 16'd-3292;
parameter WEIGHT_0_1873 = 16'd-3379;
parameter WEIGHT_0_1874 = 16'd-3978;
parameter WEIGHT_0_1875 = 16'd2048;
parameter WEIGHT_0_1876 = 16'd-651;
parameter WEIGHT_0_1877 = 16'd-6147;
parameter WEIGHT_0_1878 = 16'd770;
parameter WEIGHT_0_1879 = 16'd-1390;
parameter WEIGHT_0_1880 = 16'd4042;
parameter WEIGHT_0_1881 = 16'd-591;
parameter WEIGHT_0_1882 = 16'd-481;
parameter WEIGHT_0_1883 = 16'd180;
parameter WEIGHT_0_1884 = 16'd-2116;
parameter WEIGHT_0_1885 = 16'd2412;
parameter WEIGHT_0_1886 = 16'd-1722;
parameter WEIGHT_0_1887 = 16'd-4885;
parameter WEIGHT_0_1888 = 16'd1947;
parameter WEIGHT_0_1889 = 16'd-453;
parameter WEIGHT_0_1890 = 16'd5443;
parameter WEIGHT_0_1891 = 16'd1695;
parameter WEIGHT_0_1892 = 16'd-1489;
parameter WEIGHT_0_1893 = 16'd-3806;
parameter WEIGHT_0_1894 = 16'd1719;
parameter WEIGHT_0_1895 = 16'd3044;
parameter WEIGHT_0_1896 = 16'd-1799;
parameter WEIGHT_0_1897 = 16'd-781;
parameter WEIGHT_0_1898 = 16'd166;
parameter WEIGHT_0_1899 = 16'd-4369;
parameter WEIGHT_0_1900 = 16'd4994;
parameter WEIGHT_0_1901 = 16'd2189;
parameter WEIGHT_0_1902 = 16'd-5771;
parameter WEIGHT_0_1903 = 16'd-7971;
parameter WEIGHT_0_1904 = 16'd3171;
parameter WEIGHT_0_1905 = 16'd5256;
parameter WEIGHT_0_1906 = 16'd2900;
parameter WEIGHT_0_1907 = 16'd-6745;
parameter WEIGHT_0_1908 = 16'd-1408;
parameter WEIGHT_0_1909 = 16'd-11699;
parameter WEIGHT_0_1910 = 16'd-1658;
parameter WEIGHT_0_1911 = 16'd435;
parameter WEIGHT_0_1912 = 16'd-12544;
parameter WEIGHT_0_1913 = 16'd-10714;
parameter WEIGHT_0_1914 = 16'd11370;
parameter WEIGHT_0_1915 = 16'd5900;
parameter WEIGHT_0_1916 = 16'd1461;
parameter WEIGHT_0_1917 = 16'd-13591;
parameter WEIGHT_0_1918 = 16'd3645;
parameter WEIGHT_0_1919 = 16'd-15567;
parameter WEIGHT_0_1920 = 16'd-11895;
parameter WEIGHT_0_1921 = 16'd-4781;
parameter WEIGHT_0_1922 = 16'd-14044;
parameter WEIGHT_0_1923 = 16'd-11216;
parameter WEIGHT_0_1924 = 16'd1277;
parameter WEIGHT_0_1925 = 16'd14141;
parameter WEIGHT_0_1926 = 16'd-1121;
parameter WEIGHT_0_1927 = 16'd-17411;
parameter WEIGHT_0_1928 = 16'd-964;
parameter WEIGHT_0_1929 = 16'd-17901;
parameter WEIGHT_0_1930 = 16'd-23155;
parameter WEIGHT_0_1931 = 16'd-17881;
parameter WEIGHT_0_1932 = 16'd-12400;
parameter WEIGHT_0_1933 = 16'd-14166;
parameter WEIGHT_0_1934 = 16'd-4478;
parameter WEIGHT_0_1935 = 16'd11689;
parameter WEIGHT_0_1936 = 16'd-1348;
parameter WEIGHT_0_1937 = 16'd-17535;
parameter WEIGHT_0_1938 = 16'd1644;
parameter WEIGHT_0_1939 = 16'd-11279;
parameter WEIGHT_0_1940 = 16'd-16286;
parameter WEIGHT_0_1941 = 16'd-6483;
parameter WEIGHT_0_1942 = 16'd-11406;
parameter WEIGHT_0_1943 = 16'd-3640;
parameter WEIGHT_0_1944 = 16'd-1723;
parameter WEIGHT_0_1945 = 16'd7309;
parameter WEIGHT_0_1946 = 16'd-2767;
parameter WEIGHT_0_1947 = 16'd-8279;
parameter WEIGHT_0_1948 = 16'd-1934;
parameter WEIGHT_0_1949 = 16'd-8097;
parameter WEIGHT_0_1950 = 16'd-2487;
parameter WEIGHT_0_1951 = 16'd-4465;
parameter WEIGHT_0_1952 = 16'd-2737;
parameter WEIGHT_0_1953 = 16'd-3527;
parameter WEIGHT_0_1954 = 16'd-7520;
parameter WEIGHT_0_1955 = 16'd6857;
parameter WEIGHT_0_1956 = 16'd-2603;
parameter WEIGHT_0_1957 = 16'd-5340;
parameter WEIGHT_0_1958 = 16'd-346;
parameter WEIGHT_0_1959 = 16'd-1405;
parameter WEIGHT_0_1960 = 16'd-1577;
parameter WEIGHT_0_1961 = 16'd1240;
parameter WEIGHT_0_1962 = 16'd891;
parameter WEIGHT_0_1963 = 16'd310;
parameter WEIGHT_0_1964 = 16'd65;
parameter WEIGHT_0_1965 = 16'd-848;
parameter WEIGHT_0_1966 = 16'd-695;
parameter WEIGHT_0_1967 = 16'd2423;
parameter WEIGHT_0_1968 = 16'd-3010;
parameter WEIGHT_0_1969 = 16'd-2660;
parameter WEIGHT_0_1970 = 16'd-7719;
parameter WEIGHT_0_1971 = 16'd-2536;
parameter WEIGHT_0_1972 = 16'd-5963;
parameter WEIGHT_0_1973 = 16'd1123;
parameter WEIGHT_0_1974 = 16'd-3405;
parameter WEIGHT_0_1975 = 16'd-3673;
parameter WEIGHT_0_1976 = 16'd-2120;
parameter WEIGHT_0_1977 = 16'd4047;
parameter WEIGHT_0_1978 = 16'd-4754;
parameter WEIGHT_0_1979 = 16'd-7211;
parameter WEIGHT_0_1980 = 16'd-2604;
parameter WEIGHT_0_1981 = 16'd-2979;
parameter WEIGHT_0_1982 = 16'd3358;
parameter WEIGHT_0_1983 = 16'd-3452;
parameter WEIGHT_0_1984 = 16'd-5199;
parameter WEIGHT_0_1985 = 16'd-1479;
parameter WEIGHT_0_1986 = 16'd-2632;
parameter WEIGHT_0_1987 = 16'd7021;
parameter WEIGHT_0_1988 = 16'd-5941;
parameter WEIGHT_0_1989 = 16'd-5213;
parameter WEIGHT_0_1990 = 16'd-3561;
parameter WEIGHT_0_1991 = 16'd-3402;
parameter WEIGHT_0_1992 = 16'd2554;
parameter WEIGHT_0_1993 = 16'd4563;
parameter WEIGHT_0_1994 = 16'd-1130;
parameter WEIGHT_0_1995 = 16'd-14880;
parameter WEIGHT_0_1996 = 16'd-10316;
parameter WEIGHT_0_1997 = 16'd6923;
parameter WEIGHT_0_1998 = 16'd-11325;
parameter WEIGHT_0_1999 = 16'd-13570;
parameter WEIGHT_0_2000 = 16'd-10626;
parameter WEIGHT_0_2001 = 16'd-1880;
parameter WEIGHT_0_2002 = 16'd6185;
parameter WEIGHT_0_2003 = 16'd6614;
parameter WEIGHT_0_2004 = 16'd1882;
parameter WEIGHT_0_2005 = 16'd-17487;
parameter WEIGHT_0_2006 = 16'd-7209;
parameter WEIGHT_0_2007 = 16'd3047;
parameter WEIGHT_0_2008 = 16'd-6615;
parameter WEIGHT_0_2009 = 16'd-18170;
parameter WEIGHT_0_2010 = 16'd-4703;
parameter WEIGHT_0_2011 = 16'd-10317;
parameter WEIGHT_0_2012 = 16'd3234;
parameter WEIGHT_0_2013 = 16'd8050;
parameter WEIGHT_0_2014 = 16'd3026;
parameter WEIGHT_0_2015 = 16'd-6740;
parameter WEIGHT_0_2016 = 16'd-3527;
parameter WEIGHT_0_2017 = 16'd4284;
parameter WEIGHT_0_2018 = 16'd-6013;
parameter WEIGHT_0_2019 = 16'd-15691;
parameter WEIGHT_0_2020 = 16'd-874;
parameter WEIGHT_0_2021 = 16'd-7035;
parameter WEIGHT_0_2022 = 16'd6325;
parameter WEIGHT_0_2023 = 16'd6228;
parameter WEIGHT_0_2024 = 16'd-1149;
parameter WEIGHT_0_2025 = 16'd-3016;
parameter WEIGHT_0_2026 = 16'd-6014;
parameter WEIGHT_0_2027 = 16'd4656;
parameter WEIGHT_0_2028 = 16'd-271;
parameter WEIGHT_0_2029 = 16'd-9339;
parameter WEIGHT_0_2030 = 16'd-6022;
parameter WEIGHT_0_2031 = 16'd-9155;
parameter WEIGHT_0_2032 = 16'd1595;
parameter WEIGHT_0_2033 = 16'd520;
parameter WEIGHT_0_2034 = 16'd1095;
parameter WEIGHT_0_2035 = 16'd-1804;
parameter WEIGHT_0_2036 = 16'd-1393;
parameter WEIGHT_0_2037 = 16'd8074;
parameter WEIGHT_0_2038 = 16'd-1819;
parameter WEIGHT_0_2039 = 16'd-10528;
parameter WEIGHT_0_2040 = 16'd-8047;
parameter WEIGHT_0_2041 = 16'd-12349;
parameter WEIGHT_0_2042 = 16'd1137;
parameter WEIGHT_0_2043 = 16'd2935;
parameter WEIGHT_0_2044 = 16'd-2187;
parameter WEIGHT_0_2045 = 16'd2560;
parameter WEIGHT_0_2046 = 16'd-3436;
parameter WEIGHT_0_2047 = 16'd5761;
parameter WEIGHT_0_2048 = 16'd1977;
parameter WEIGHT_0_2049 = 16'd-3004;
parameter WEIGHT_0_2050 = 16'd-2895;
parameter WEIGHT_0_2051 = 16'd-8450;
parameter WEIGHT_0_2052 = 16'd1013;
parameter WEIGHT_0_2053 = 16'd1184;
parameter WEIGHT_0_2054 = 16'd-2738;
parameter WEIGHT_0_2055 = 16'd3607;
parameter WEIGHT_0_2056 = 16'd-3832;
parameter WEIGHT_0_2057 = 16'd4169;
parameter WEIGHT_0_2058 = 16'd-461;
parameter WEIGHT_0_2059 = 16'd-5119;
parameter WEIGHT_0_2060 = 16'd-874;
parameter WEIGHT_0_2061 = 16'd-6931;
parameter WEIGHT_0_2062 = 16'd1110;
parameter WEIGHT_0_2063 = 16'd3047;
parameter WEIGHT_0_2064 = 16'd-5482;
parameter WEIGHT_0_2065 = 16'd2859;
parameter WEIGHT_0_2066 = 16'd-3173;
parameter WEIGHT_0_2067 = 16'd4550;
parameter WEIGHT_0_2068 = 16'd362;
parameter WEIGHT_0_2069 = 16'd-868;
parameter WEIGHT_0_2070 = 16'd-1736;
parameter WEIGHT_0_2071 = 16'd-4531;
parameter WEIGHT_0_2072 = 16'd2447;
parameter WEIGHT_0_2073 = 16'd3077;
parameter WEIGHT_0_2074 = 16'd-7891;
parameter WEIGHT_0_2075 = 16'd6696;
parameter WEIGHT_0_2076 = 16'd-2632;
parameter WEIGHT_0_2077 = 16'd7452;
parameter WEIGHT_0_2078 = 16'd326;
parameter WEIGHT_0_2079 = 16'd119;
parameter WEIGHT_0_2080 = 16'd2836;
parameter WEIGHT_0_2081 = 16'd-3692;
parameter WEIGHT_0_2082 = 16'd1026;
parameter WEIGHT_0_2083 = 16'd5123;
parameter WEIGHT_0_2084 = 16'd-9924;
parameter WEIGHT_0_2085 = 16'd1124;
parameter WEIGHT_0_2086 = 16'd-3376;
parameter WEIGHT_0_2087 = 16'd3252;
parameter WEIGHT_0_2088 = 16'd-172;
parameter WEIGHT_0_2089 = 16'd2283;
parameter WEIGHT_0_2090 = 16'd3168;
parameter WEIGHT_0_2091 = 16'd-3256;
parameter WEIGHT_0_2092 = 16'd196;
parameter WEIGHT_0_2093 = 16'd3203;
parameter WEIGHT_0_2094 = 16'd-8627;
parameter WEIGHT_0_2095 = 16'd-395;
parameter WEIGHT_0_2096 = 16'd-4036;
parameter WEIGHT_0_2097 = 16'd3999;
parameter WEIGHT_0_2098 = 16'd-1068;
parameter WEIGHT_0_2099 = 16'd8325;
parameter WEIGHT_0_2100 = 16'd811;
parameter WEIGHT_0_2101 = 16'd-2649;
parameter WEIGHT_0_2102 = 16'd3560;
parameter WEIGHT_0_2103 = 16'd3950;
parameter WEIGHT_0_2104 = 16'd-14512;
parameter WEIGHT_0_2105 = 16'd117;
parameter WEIGHT_0_2106 = 16'd-6059;
parameter WEIGHT_0_2107 = 16'd-1885;
parameter WEIGHT_0_2108 = 16'd-3034;
parameter WEIGHT_0_2109 = 16'd10124;
parameter WEIGHT_0_2110 = 16'd4067;
parameter WEIGHT_0_2111 = 16'd-6819;
parameter WEIGHT_0_2112 = 16'd-2914;
parameter WEIGHT_0_2113 = 16'd4798;
parameter WEIGHT_0_2114 = 16'd-14327;
parameter WEIGHT_0_2115 = 16'd-1781;
parameter WEIGHT_0_2116 = 16'd-7102;
parameter WEIGHT_0_2117 = 16'd-340;
parameter WEIGHT_0_2118 = 16'd508;
parameter WEIGHT_0_2119 = 16'd14052;
parameter WEIGHT_0_2120 = 16'd5376;
parameter WEIGHT_0_2121 = 16'd-7111;
parameter WEIGHT_0_2122 = 16'd2017;
parameter WEIGHT_0_2123 = 16'd1016;
parameter WEIGHT_0_2124 = 16'd-11405;
parameter WEIGHT_0_2125 = 16'd-341;
parameter WEIGHT_0_2126 = 16'd-5839;
parameter WEIGHT_0_2127 = 16'd1858;
parameter WEIGHT_0_2128 = 16'd2409;
parameter WEIGHT_0_2129 = 16'd10881;
parameter WEIGHT_0_2130 = 16'd8091;
parameter WEIGHT_0_2131 = 16'd-4599;
parameter WEIGHT_0_2132 = 16'd-5030;
parameter WEIGHT_0_2133 = 16'd4229;
parameter WEIGHT_0_2134 = 16'd-8408;
parameter WEIGHT_0_2135 = 16'd2032;
parameter WEIGHT_0_2136 = 16'd-9487;
parameter WEIGHT_0_2137 = 16'd3937;
parameter WEIGHT_0_2138 = 16'd-387;
parameter WEIGHT_0_2139 = 16'd4426;
parameter WEIGHT_0_2140 = 16'd7594;
parameter WEIGHT_0_2141 = 16'd-5324;
parameter WEIGHT_0_2142 = 16'd-217;
parameter WEIGHT_0_2143 = 16'd3590;
parameter WEIGHT_0_2144 = 16'd-8955;
parameter WEIGHT_0_2145 = 16'd3328;
parameter WEIGHT_0_2146 = 16'd-8390;
parameter WEIGHT_0_2147 = 16'd6697;
parameter WEIGHT_0_2148 = 16'd-231;
parameter WEIGHT_0_2149 = 16'd3138;
parameter WEIGHT_0_2150 = 16'd2718;
parameter WEIGHT_0_2151 = 16'd-661;
parameter WEIGHT_0_2152 = 16'd-2705;
parameter WEIGHT_0_2153 = 16'd-982;
parameter WEIGHT_0_2154 = 16'd-5222;
parameter WEIGHT_0_2155 = 16'd1291;
parameter WEIGHT_0_2156 = 16'd-6959;
parameter WEIGHT_0_2157 = 16'd777;
parameter WEIGHT_0_2158 = 16'd-900;
parameter WEIGHT_0_2159 = 16'd-1037;
parameter WEIGHT_0_2160 = 16'd161;
parameter WEIGHT_0_2161 = 16'd771;
parameter WEIGHT_0_2162 = 16'd-2945;
parameter WEIGHT_0_2163 = 16'd2215;
parameter WEIGHT_0_2164 = 16'd-2968;
parameter WEIGHT_0_2165 = 16'd3558;
parameter WEIGHT_0_2166 = 16'd-5926;
parameter WEIGHT_0_2167 = 16'd2246;
parameter WEIGHT_0_2168 = 16'd1743;
parameter WEIGHT_0_2169 = 16'd-1658;
parameter WEIGHT_0_2170 = 16'd-304;
parameter WEIGHT_0_2171 = 16'd-2676;
parameter WEIGHT_0_2172 = 16'd969;
parameter WEIGHT_0_2173 = 16'd-2433;
parameter WEIGHT_0_2174 = 16'd-1685;
parameter WEIGHT_0_2175 = 16'd2651;
parameter WEIGHT_0_2176 = 16'd-2434;
parameter WEIGHT_0_2177 = 16'd-538;
parameter WEIGHT_0_2178 = 16'd4024;
parameter WEIGHT_0_2179 = 16'd-3309;
parameter WEIGHT_0_2180 = 16'd4235;
parameter WEIGHT_0_2181 = 16'd-4508;
parameter WEIGHT_0_2182 = 16'd2273;
parameter WEIGHT_0_2183 = 16'd-4345;
parameter WEIGHT_0_2184 = 16'd5144;
parameter WEIGHT_0_2185 = 16'd6163;
parameter WEIGHT_0_2186 = 16'd-6666;
parameter WEIGHT_0_2187 = 16'd-2535;
parameter WEIGHT_0_2188 = 16'd2525;
parameter WEIGHT_0_2189 = 16'd-7096;
parameter WEIGHT_0_2190 = 16'd889;
parameter WEIGHT_0_2191 = 16'd-3632;
parameter WEIGHT_0_2192 = 16'd-11956;
parameter WEIGHT_0_2193 = 16'd-12680;
parameter WEIGHT_0_2194 = 16'd6148;
parameter WEIGHT_0_2195 = 16'd8920;
parameter WEIGHT_0_2196 = 16'd-4775;
parameter WEIGHT_0_2197 = 16'd-4087;
parameter WEIGHT_0_2198 = 16'd2527;
parameter WEIGHT_0_2199 = 16'd-15219;
parameter WEIGHT_0_2200 = 16'd-7238;
parameter WEIGHT_0_2201 = 16'd-16081;
parameter WEIGHT_0_2202 = 16'd-21382;
parameter WEIGHT_0_2203 = 16'd-16507;
parameter WEIGHT_0_2204 = 16'd1613;
parameter WEIGHT_0_2205 = 16'd14602;
parameter WEIGHT_0_2206 = 16'd-4706;
parameter WEIGHT_0_2207 = 16'd-11745;
parameter WEIGHT_0_2208 = 16'd2979;
parameter WEIGHT_0_2209 = 16'd-16258;
parameter WEIGHT_0_2210 = 16'd-23040;
parameter WEIGHT_0_2211 = 16'd-21767;
parameter WEIGHT_0_2212 = 16'd-10173;
parameter WEIGHT_0_2213 = 16'd-20938;
parameter WEIGHT_0_2214 = 16'd-3277;
parameter WEIGHT_0_2215 = 16'd15579;
parameter WEIGHT_0_2216 = 16'd-3244;
parameter WEIGHT_0_2217 = 16'd-13346;
parameter WEIGHT_0_2218 = 16'd-3904;
parameter WEIGHT_0_2219 = 16'd-14931;
parameter WEIGHT_0_2220 = 16'd-17237;
parameter WEIGHT_0_2221 = 16'd-9806;
parameter WEIGHT_0_2222 = 16'd-8506;
parameter WEIGHT_0_2223 = 16'd-6429;
parameter WEIGHT_0_2224 = 16'd-332;
parameter WEIGHT_0_2225 = 16'd7562;
parameter WEIGHT_0_2226 = 16'd-5482;
parameter WEIGHT_0_2227 = 16'd-8009;
parameter WEIGHT_0_2228 = 16'd-300;
parameter WEIGHT_0_2229 = 16'd-13463;
parameter WEIGHT_0_2230 = 16'd-1904;
parameter WEIGHT_0_2231 = 16'd-2527;
parameter WEIGHT_0_2232 = 16'd-7024;
parameter WEIGHT_0_2233 = 16'd301;
parameter WEIGHT_0_2234 = 16'd-5361;
parameter WEIGHT_0_2235 = 16'd4102;
parameter WEIGHT_0_2236 = 16'd-1887;
parameter WEIGHT_0_2237 = 16'd-6142;
parameter WEIGHT_0_2238 = 16'd46;
parameter WEIGHT_0_2239 = 16'd-6365;
parameter WEIGHT_0_2240 = 16'd723;
parameter WEIGHT_0_2241 = 16'd-3119;
parameter WEIGHT_0_2242 = 16'd-803;
parameter WEIGHT_0_2243 = 16'd-2469;
parameter WEIGHT_0_2244 = 16'd-3924;
parameter WEIGHT_0_2245 = 16'd-2707;
parameter WEIGHT_0_2246 = 16'd-815;
parameter WEIGHT_0_2247 = 16'd-1765;
parameter WEIGHT_0_2248 = 16'd-1843;
parameter WEIGHT_0_2249 = 16'd-4927;
parameter WEIGHT_0_2250 = 16'd-6518;
parameter WEIGHT_0_2251 = 16'd-4440;
parameter WEIGHT_0_2252 = 16'd1173;
parameter WEIGHT_0_2253 = 16'd-4758;
parameter WEIGHT_0_2254 = 16'd-6473;
parameter WEIGHT_0_2255 = 16'd-5876;
parameter WEIGHT_0_2256 = 16'd915;
parameter WEIGHT_0_2257 = 16'd3600;
parameter WEIGHT_0_2258 = 16'd-4024;
parameter WEIGHT_0_2259 = 16'd-3754;
parameter WEIGHT_0_2260 = 16'd-723;
parameter WEIGHT_0_2261 = 16'd-1693;
parameter WEIGHT_0_2262 = 16'd-949;
parameter WEIGHT_0_2263 = 16'd-4442;
parameter WEIGHT_0_2264 = 16'd567;
parameter WEIGHT_0_2265 = 16'd-6914;
parameter WEIGHT_0_2266 = 16'd-4396;
parameter WEIGHT_0_2267 = 16'd7213;
parameter WEIGHT_0_2268 = 16'd-6560;
parameter WEIGHT_0_2269 = 16'd-11957;
parameter WEIGHT_0_2270 = 16'd-4265;
parameter WEIGHT_0_2271 = 16'd-184;
parameter WEIGHT_0_2272 = 16'd-333;
parameter WEIGHT_0_2273 = 16'd3423;
parameter WEIGHT_0_2274 = 16'd-1963;
parameter WEIGHT_0_2275 = 16'd-16940;
parameter WEIGHT_0_2276 = 16'd-7837;
parameter WEIGHT_0_2277 = 16'd8689;
parameter WEIGHT_0_2278 = 16'd-1636;
parameter WEIGHT_0_2279 = 16'd-13964;
parameter WEIGHT_0_2280 = 16'd-12270;
parameter WEIGHT_0_2281 = 16'd-3475;
parameter WEIGHT_0_2282 = 16'd4173;
parameter WEIGHT_0_2283 = 16'd8565;
parameter WEIGHT_0_2284 = 16'd-1337;
parameter WEIGHT_0_2285 = 16'd-18164;
parameter WEIGHT_0_2286 = 16'd-1249;
parameter WEIGHT_0_2287 = 16'd4021;
parameter WEIGHT_0_2288 = 16'd-4265;
parameter WEIGHT_0_2289 = 16'd-14828;
parameter WEIGHT_0_2290 = 16'd-7194;
parameter WEIGHT_0_2291 = 16'd-7702;
parameter WEIGHT_0_2292 = 16'd2025;
parameter WEIGHT_0_2293 = 16'd4995;
parameter WEIGHT_0_2294 = 16'd-279;
parameter WEIGHT_0_2295 = 16'd-9620;
parameter WEIGHT_0_2296 = 16'd-5477;
parameter WEIGHT_0_2297 = 16'd5452;
parameter WEIGHT_0_2298 = 16'd-2598;
parameter WEIGHT_0_2299 = 16'd-9415;
parameter WEIGHT_0_2300 = 16'd-3230;
parameter WEIGHT_0_2301 = 16'd-8419;
parameter WEIGHT_0_2302 = 16'd629;
parameter WEIGHT_0_2303 = 16'd3570;
parameter WEIGHT_0_2304 = 16'd-1926;
parameter WEIGHT_0_2305 = 16'd-3956;
parameter WEIGHT_0_2306 = 16'd-8313;
parameter WEIGHT_0_2307 = 16'd4333;
parameter WEIGHT_0_2308 = 16'd1660;
parameter WEIGHT_0_2309 = 16'd-6278;
parameter WEIGHT_0_2310 = 16'd-3877;
parameter WEIGHT_0_2311 = 16'd-6584;
parameter WEIGHT_0_2312 = 16'd1968;
parameter WEIGHT_0_2313 = 16'd2560;
parameter WEIGHT_0_2314 = 16'd-1687;
parameter WEIGHT_0_2315 = 16'd-3427;
parameter WEIGHT_0_2316 = 16'd-1375;
parameter WEIGHT_0_2317 = 16'd5979;
parameter WEIGHT_0_2318 = 16'd2144;
parameter WEIGHT_0_2319 = 16'd-7320;
parameter WEIGHT_0_2320 = 16'd-961;
parameter WEIGHT_0_2321 = 16'd-11156;
parameter WEIGHT_0_2322 = 16'd2657;
parameter WEIGHT_0_2323 = 16'd-1425;
parameter WEIGHT_0_2324 = 16'd-5218;
parameter WEIGHT_0_2325 = 16'd3227;
parameter WEIGHT_0_2326 = 16'd-4455;
parameter WEIGHT_0_2327 = 16'd7385;
parameter WEIGHT_0_2328 = 16'd862;
parameter WEIGHT_0_2329 = 16'd-1239;
parameter WEIGHT_0_2330 = 16'd1962;
parameter WEIGHT_0_2331 = 16'd-11491;
parameter WEIGHT_0_2332 = 16'd1282;
parameter WEIGHT_0_2333 = 16'd1666;
parameter WEIGHT_0_2334 = 16'd-3157;
parameter WEIGHT_0_2335 = 16'd2835;
parameter WEIGHT_0_2336 = 16'd-3199;
parameter WEIGHT_0_2337 = 16'd6306;
parameter WEIGHT_0_2338 = 16'd1515;
parameter WEIGHT_0_2339 = 16'd-2976;
parameter WEIGHT_0_2340 = 16'd-1836;
parameter WEIGHT_0_2341 = 16'd-9037;
parameter WEIGHT_0_2342 = 16'd5457;
parameter WEIGHT_0_2343 = 16'd-2155;
parameter WEIGHT_0_2344 = 16'd-3359;
parameter WEIGHT_0_2345 = 16'd1587;
parameter WEIGHT_0_2346 = 16'd-7109;
parameter WEIGHT_0_2347 = 16'd5945;
parameter WEIGHT_0_2348 = 16'd3874;
parameter WEIGHT_0_2349 = 16'd-845;
parameter WEIGHT_0_2350 = 16'd539;
parameter WEIGHT_0_2351 = 16'd-5858;
parameter WEIGHT_0_2352 = 16'd4352;
parameter WEIGHT_0_2353 = 16'd-1075;
parameter WEIGHT_0_2354 = 16'd-5450;
parameter WEIGHT_0_2355 = 16'd1976;
parameter WEIGHT_0_2356 = 16'd-4744;
parameter WEIGHT_0_2357 = 16'd6959;
parameter WEIGHT_0_2358 = 16'd-301;
parameter WEIGHT_0_2359 = 16'd-3981;
parameter WEIGHT_0_2360 = 16'd-599;
parameter WEIGHT_0_2361 = 16'd-2167;
parameter WEIGHT_0_2362 = 16'd1567;
parameter WEIGHT_0_2363 = 16'd757;
parameter WEIGHT_0_2364 = 16'd-7579;
parameter WEIGHT_0_2365 = 16'd472;
parameter WEIGHT_0_2366 = 16'd-3957;
parameter WEIGHT_0_2367 = 16'd7769;
parameter WEIGHT_0_2368 = 16'd3735;
parameter WEIGHT_0_2369 = 16'd147;
parameter WEIGHT_0_2370 = 16'd1231;
parameter WEIGHT_0_2371 = 16'd-407;
parameter WEIGHT_0_2372 = 16'd1114;
parameter WEIGHT_0_2373 = 16'd1933;
parameter WEIGHT_0_2374 = 16'd-6924;
parameter WEIGHT_0_2375 = 16'd449;
parameter WEIGHT_0_2376 = 16'd-5004;
parameter WEIGHT_0_2377 = 16'd2733;
parameter WEIGHT_0_2378 = 16'd3061;
parameter WEIGHT_0_2379 = 16'd4575;
parameter WEIGHT_0_2380 = 16'd3714;
parameter WEIGHT_0_2381 = 16'd-2498;
parameter WEIGHT_0_2382 = 16'd3072;
parameter WEIGHT_0_2383 = 16'd4794;
parameter WEIGHT_0_2384 = 16'd-14696;
parameter WEIGHT_0_2385 = 16'd-3917;
parameter WEIGHT_0_2386 = 16'd-4754;
parameter WEIGHT_0_2387 = 16'd4925;
parameter WEIGHT_0_2388 = 16'd-3031;
parameter WEIGHT_0_2389 = 16'd4475;
parameter WEIGHT_0_2390 = 16'd5002;
parameter WEIGHT_0_2391 = 16'd1460;
parameter WEIGHT_0_2392 = 16'd4215;
parameter WEIGHT_0_2393 = 16'd4079;
parameter WEIGHT_0_2394 = 16'd-14353;
parameter WEIGHT_0_2395 = 16'd-7221;
parameter WEIGHT_0_2396 = 16'd-6995;
parameter WEIGHT_0_2397 = 16'd4471;
parameter WEIGHT_0_2398 = 16'd-2109;
parameter WEIGHT_0_2399 = 16'd7650;
parameter WEIGHT_0_2400 = 16'd5896;
parameter WEIGHT_0_2401 = 16'd-2990;
parameter WEIGHT_0_2402 = 16'd524;
parameter WEIGHT_0_2403 = 16'd5536;
parameter WEIGHT_0_2404 = 16'd-11106;
parameter WEIGHT_0_2405 = 16'd-3112;
parameter WEIGHT_0_2406 = 16'd-7515;
parameter WEIGHT_0_2407 = 16'd8849;
parameter WEIGHT_0_2408 = 16'd-2210;
parameter WEIGHT_0_2409 = 16'd5700;
parameter WEIGHT_0_2410 = 16'd8307;
parameter WEIGHT_0_2411 = 16'd-1019;
parameter WEIGHT_0_2412 = 16'd-515;
parameter WEIGHT_0_2413 = 16'd1849;
parameter WEIGHT_0_2414 = 16'd-5735;
parameter WEIGHT_0_2415 = 16'd-3370;
parameter WEIGHT_0_2416 = 16'd-12658;
parameter WEIGHT_0_2417 = 16'd8495;
parameter WEIGHT_0_2418 = 16'd-719;
parameter WEIGHT_0_2419 = 16'd2408;
parameter WEIGHT_0_2420 = 16'd7245;
parameter WEIGHT_0_2421 = 16'd-2558;
parameter WEIGHT_0_2422 = 16'd-2849;
parameter WEIGHT_0_2423 = 16'd2897;
parameter WEIGHT_0_2424 = 16'd-2521;
parameter WEIGHT_0_2425 = 16'd-2914;
parameter WEIGHT_0_2426 = 16'd-13860;
parameter WEIGHT_0_2427 = 16'd5947;
parameter WEIGHT_0_2428 = 16'd2239;
parameter WEIGHT_0_2429 = 16'd1426;
parameter WEIGHT_0_2430 = 16'd4245;
parameter WEIGHT_0_2431 = 16'd-1938;
parameter WEIGHT_0_2432 = 16'd2234;
parameter WEIGHT_0_2433 = 16'd1268;
parameter WEIGHT_0_2434 = 16'd-3790;
parameter WEIGHT_0_2435 = 16'd1544;
parameter WEIGHT_0_2436 = 16'd-15277;
parameter WEIGHT_0_2437 = 16'd2643;
parameter WEIGHT_0_2438 = 16'd3259;
parameter WEIGHT_0_2439 = 16'd-4531;
parameter WEIGHT_0_2440 = 16'd3036;
parameter WEIGHT_0_2441 = 16'd-3677;
parameter WEIGHT_0_2442 = 16'd-2152;
parameter WEIGHT_0_2443 = 16'd1947;
parameter WEIGHT_0_2444 = 16'd-1008;
parameter WEIGHT_0_2445 = 16'd4070;
parameter WEIGHT_0_2446 = 16'd-9514;
parameter WEIGHT_0_2447 = 16'd1853;
parameter WEIGHT_0_2448 = 16'd783;
parameter WEIGHT_0_2449 = 16'd-4353;
parameter WEIGHT_0_2450 = 16'd2910;
parameter WEIGHT_0_2451 = 16'd-3562;
parameter WEIGHT_0_2452 = 16'd-2661;
parameter WEIGHT_0_2453 = 16'd-1741;
parameter WEIGHT_0_2454 = 16'd-1170;
parameter WEIGHT_0_2455 = 16'd7014;
parameter WEIGHT_0_2456 = 16'd-7050;
parameter WEIGHT_0_2457 = 16'd-2451;
parameter WEIGHT_0_2458 = 16'd2270;
parameter WEIGHT_0_2459 = 16'd-854;
parameter WEIGHT_0_2460 = 16'd3682;
parameter WEIGHT_0_2461 = 16'd-7277;
parameter WEIGHT_0_2462 = 16'd-2340;
parameter WEIGHT_0_2463 = 16'd2476;
parameter WEIGHT_0_2464 = 16'd-129;
parameter WEIGHT_0_2465 = 16'd4308;
parameter WEIGHT_0_2466 = 16'd-8433;
parameter WEIGHT_0_2467 = 16'd1222;
parameter WEIGHT_0_2468 = 16'd6243;
parameter WEIGHT_0_2469 = 16'd-5605;
parameter WEIGHT_0_2470 = 16'd3794;
parameter WEIGHT_0_2471 = 16'd-14341;
parameter WEIGHT_0_2472 = 16'd-5172;
parameter WEIGHT_0_2473 = 16'd-11456;
parameter WEIGHT_0_2474 = 16'd1195;
parameter WEIGHT_0_2475 = 16'd11090;
parameter WEIGHT_0_2476 = 16'd-10733;
parameter WEIGHT_0_2477 = 16'd-4155;
parameter WEIGHT_0_2478 = 16'd4922;
parameter WEIGHT_0_2479 = 16'd-9347;
parameter WEIGHT_0_2480 = 16'd-876;
parameter WEIGHT_0_2481 = 16'd-20119;
parameter WEIGHT_0_2482 = 16'd-22870;
parameter WEIGHT_0_2483 = 16'd-28680;
parameter WEIGHT_0_2484 = 16'd-4772;
parameter WEIGHT_0_2485 = 16'd21234;
parameter WEIGHT_0_2486 = 16'd-13772;
parameter WEIGHT_0_2487 = 16'd-12935;
parameter WEIGHT_0_2488 = 16'd3925;
parameter WEIGHT_0_2489 = 16'd-13420;
parameter WEIGHT_0_2490 = 16'd-22370;
parameter WEIGHT_0_2491 = 16'd-22222;
parameter WEIGHT_0_2492 = 16'd-21797;
parameter WEIGHT_0_2493 = 16'd-21604;
parameter WEIGHT_0_2494 = 16'd-3258;
parameter WEIGHT_0_2495 = 16'd19737;
parameter WEIGHT_0_2496 = 16'd-16162;
parameter WEIGHT_0_2497 = 16'd-16548;
parameter WEIGHT_0_2498 = 16'd1273;
parameter WEIGHT_0_2499 = 16'd-13806;
parameter WEIGHT_0_2500 = 16'd-14616;
parameter WEIGHT_0_2501 = 16'd-7146;
parameter WEIGHT_0_2502 = 16'd-10495;
parameter WEIGHT_0_2503 = 16'd-9124;
parameter WEIGHT_0_2504 = 16'd-1981;
parameter WEIGHT_0_2505 = 16'd11215;
parameter WEIGHT_0_2506 = 16'd-12270;
parameter WEIGHT_0_2507 = 16'd-9386;
parameter WEIGHT_0_2508 = 16'd3046;
parameter WEIGHT_0_2509 = 16'd-11912;
parameter WEIGHT_0_2510 = 16'd-4652;
parameter WEIGHT_0_2511 = 16'd-1011;
parameter WEIGHT_0_2512 = 16'd-6178;
parameter WEIGHT_0_2513 = 16'd-2615;
parameter WEIGHT_0_2514 = 16'd-3083;
parameter WEIGHT_0_2515 = 16'd4093;
parameter WEIGHT_0_2516 = 16'd-6265;
parameter WEIGHT_0_2517 = 16'd-1286;
parameter WEIGHT_0_2518 = 16'd1052;
parameter WEIGHT_0_2519 = 16'd-2876;
parameter WEIGHT_0_2520 = 16'd-4024;
parameter WEIGHT_0_2521 = 16'd-1485;
parameter WEIGHT_0_2522 = 16'd-1255;
parameter WEIGHT_0_2523 = 16'd-2387;
parameter WEIGHT_0_2524 = 16'd-4934;
parameter WEIGHT_0_2525 = 16'd-3726;
parameter WEIGHT_0_2526 = 16'd-774;
parameter WEIGHT_0_2527 = 16'd1689;
parameter WEIGHT_0_2528 = 16'd-2426;
parameter WEIGHT_0_2529 = 16'd-3493;
parameter WEIGHT_0_2530 = 16'd203;
parameter WEIGHT_0_2531 = 16'd362;
parameter WEIGHT_0_2532 = 16'd-1848;
parameter WEIGHT_0_2533 = 16'd-2617;
parameter WEIGHT_0_2534 = 16'd-2214;
parameter WEIGHT_0_2535 = 16'd-5587;
parameter WEIGHT_0_2536 = 16'd1348;
parameter WEIGHT_0_2537 = 16'd5494;
parameter WEIGHT_0_2538 = 16'd-3649;
parameter WEIGHT_0_2539 = 16'd-4965;
parameter WEIGHT_0_2540 = 16'd3802;
parameter WEIGHT_0_2541 = 16'd-1326;
parameter WEIGHT_0_2542 = 16'd-1048;
parameter WEIGHT_0_2543 = 16'd79;
parameter WEIGHT_0_2544 = 16'd-2437;
parameter WEIGHT_0_2545 = 16'd-6954;
parameter WEIGHT_0_2546 = 16'd-2466;
parameter WEIGHT_0_2547 = 16'd6676;
parameter WEIGHT_0_2548 = 16'd-8138;
parameter WEIGHT_0_2549 = 16'd-8963;
parameter WEIGHT_0_2550 = 16'd-1412;
parameter WEIGHT_0_2551 = 16'd-5934;
parameter WEIGHT_0_2552 = 16'd1378;
parameter WEIGHT_0_2553 = 16'd4373;
parameter WEIGHT_0_2554 = 16'd-10503;
parameter WEIGHT_0_2555 = 16'd-16085;
parameter WEIGHT_0_2556 = 16'd-8144;
parameter WEIGHT_0_2557 = 16'd8909;
parameter WEIGHT_0_2558 = 16'd-1951;
parameter WEIGHT_0_2559 = 16'd-8785;
parameter WEIGHT_0_2560 = 16'd-6344;
parameter WEIGHT_0_2561 = 16'd-2605;
parameter WEIGHT_0_2562 = 16'd6488;
parameter WEIGHT_0_2563 = 16'd10705;
parameter WEIGHT_0_2564 = 16'd-6204;
parameter WEIGHT_0_2565 = 16'd-14953;
parameter WEIGHT_0_2566 = 16'd-1789;
parameter WEIGHT_0_2567 = 16'd8161;
parameter WEIGHT_0_2568 = 16'd116;
parameter WEIGHT_0_2569 = 16'd-10549;
parameter WEIGHT_0_2570 = 16'd-2118;
parameter WEIGHT_0_2571 = 16'd-8194;
parameter WEIGHT_0_2572 = 16'd5428;
parameter WEIGHT_0_2573 = 16'd4358;
parameter WEIGHT_0_2574 = 16'd-3151;
parameter WEIGHT_0_2575 = 16'd-9212;
parameter WEIGHT_0_2576 = 16'd-9532;
parameter WEIGHT_0_2577 = 16'd5519;
parameter WEIGHT_0_2578 = 16'd3046;
parameter WEIGHT_0_2579 = 16'd-6099;
parameter WEIGHT_0_2580 = 16'd-3779;
parameter WEIGHT_0_2581 = 16'd-6035;
parameter WEIGHT_0_2582 = 16'd781;
parameter WEIGHT_0_2583 = 16'd3901;
parameter WEIGHT_0_2584 = 16'd-5166;
parameter WEIGHT_0_2585 = 16'd-2009;
parameter WEIGHT_0_2586 = 16'd-6378;
parameter WEIGHT_0_2587 = 16'd5449;
parameter WEIGHT_0_2588 = 16'd1157;
parameter WEIGHT_0_2589 = 16'd342;
parameter WEIGHT_0_2590 = 16'd-2805;
parameter WEIGHT_0_2591 = 16'd-3697;
parameter WEIGHT_0_2592 = 16'd-2971;
parameter WEIGHT_0_2593 = 16'd2298;
parameter WEIGHT_0_2594 = 16'd-2360;
parameter WEIGHT_0_2595 = 16'd-2121;
parameter WEIGHT_0_2596 = 16'd-2375;
parameter WEIGHT_0_2597 = 16'd1324;
parameter WEIGHT_0_2598 = 16'd5563;
parameter WEIGHT_0_2599 = 16'd-1612;
parameter WEIGHT_0_2600 = 16'd-4839;
parameter WEIGHT_0_2601 = 16'd-6032;
parameter WEIGHT_0_2602 = 16'd-618;
parameter WEIGHT_0_2603 = 16'd-2273;
parameter WEIGHT_0_2604 = 16'd-1337;
parameter WEIGHT_0_2605 = 16'd2065;
parameter WEIGHT_0_2606 = 16'd-2023;
parameter WEIGHT_0_2607 = 16'd164;
parameter WEIGHT_0_2608 = 16'd4307;
parameter WEIGHT_0_2609 = 16'd-62;
parameter WEIGHT_0_2610 = 16'd-119;
parameter WEIGHT_0_2611 = 16'd-7381;
parameter WEIGHT_0_2612 = 16'd-574;
parameter WEIGHT_0_2613 = 16'd-2086;
parameter WEIGHT_0_2614 = 16'd-711;
parameter WEIGHT_0_2615 = 16'd551;
parameter WEIGHT_0_2616 = 16'd-6715;
parameter WEIGHT_0_2617 = 16'd-1094;
parameter WEIGHT_0_2618 = 16'd5268;
parameter WEIGHT_0_2619 = 16'd-3528;
parameter WEIGHT_0_2620 = 16'd1605;
parameter WEIGHT_0_2621 = 16'd-5107;
parameter WEIGHT_0_2622 = 16'd3369;
parameter WEIGHT_0_2623 = 16'd-5334;
parameter WEIGHT_0_2624 = 16'd-3775;
parameter WEIGHT_0_2625 = 16'd4762;
parameter WEIGHT_0_2626 = 16'd-2953;
parameter WEIGHT_0_2627 = 16'd683;
parameter WEIGHT_0_2628 = 16'd2203;
parameter WEIGHT_0_2629 = 16'd-128;
parameter WEIGHT_0_2630 = 16'd-2918;
parameter WEIGHT_0_2631 = 16'd-4047;
parameter WEIGHT_0_2632 = 16'd-230;
parameter WEIGHT_0_2633 = 16'd-10135;
parameter WEIGHT_0_2634 = 16'd-3106;
parameter WEIGHT_0_2635 = 16'd8531;
parameter WEIGHT_0_2636 = 16'd-5772;
parameter WEIGHT_0_2637 = 16'd1974;
parameter WEIGHT_0_2638 = 16'd4350;
parameter WEIGHT_0_2639 = 16'd-1147;
parameter WEIGHT_0_2640 = 16'd1752;
parameter WEIGHT_0_2641 = 16'd-4109;
parameter WEIGHT_0_2642 = 16'd-223;
parameter WEIGHT_0_2643 = 16'd-6277;
parameter WEIGHT_0_2644 = 16'd-3358;
parameter WEIGHT_0_2645 = 16'd4909;
parameter WEIGHT_0_2646 = 16'd-5894;
parameter WEIGHT_0_2647 = 16'd4551;
parameter WEIGHT_0_2648 = 16'd-1278;
parameter WEIGHT_0_2649 = 16'd-2324;
parameter WEIGHT_0_2650 = 16'd4275;
parameter WEIGHT_0_2651 = 16'd3245;
parameter WEIGHT_0_2652 = 16'd609;
parameter WEIGHT_0_2653 = 16'd-1665;
parameter WEIGHT_0_2654 = 16'd-4009;
parameter WEIGHT_0_2655 = 16'd1134;
parameter WEIGHT_0_2656 = 16'd-6253;
parameter WEIGHT_0_2657 = 16'd1994;
parameter WEIGHT_0_2658 = 16'd1513;
parameter WEIGHT_0_2659 = 16'd2289;
parameter WEIGHT_0_2660 = 16'd-301;
parameter WEIGHT_0_2661 = 16'd7275;
parameter WEIGHT_0_2662 = 16'd2411;
parameter WEIGHT_0_2663 = 16'd3382;
parameter WEIGHT_0_2664 = 16'd-15125;
parameter WEIGHT_0_2665 = 16'd-5787;
parameter WEIGHT_0_2666 = 16'd-5792;
parameter WEIGHT_0_2667 = 16'd8371;
parameter WEIGHT_0_2668 = 16'd-6775;
parameter WEIGHT_0_2669 = 16'd1567;
parameter WEIGHT_0_2670 = 16'd1321;
parameter WEIGHT_0_2671 = 16'd10323;
parameter WEIGHT_0_2672 = 16'd1726;
parameter WEIGHT_0_2673 = 16'd9943;
parameter WEIGHT_0_2674 = 16'd-12093;
parameter WEIGHT_0_2675 = 16'd-7169;
parameter WEIGHT_0_2676 = 16'd-12569;
parameter WEIGHT_0_2677 = 16'd8547;
parameter WEIGHT_0_2678 = 16'd-10438;
parameter WEIGHT_0_2679 = 16'd847;
parameter WEIGHT_0_2680 = 16'd2686;
parameter WEIGHT_0_2681 = 16'd4791;
parameter WEIGHT_0_2682 = 16'd1248;
parameter WEIGHT_0_2683 = 16'd3444;
parameter WEIGHT_0_2684 = 16'd-6864;
parameter WEIGHT_0_2685 = 16'd-8721;
parameter WEIGHT_0_2686 = 16'd-11685;
parameter WEIGHT_0_2687 = 16'd8062;
parameter WEIGHT_0_2688 = 16'd-4884;
parameter WEIGHT_0_2689 = 16'd-3459;
parameter WEIGHT_0_2690 = 16'd6503;
parameter WEIGHT_0_2691 = 16'd454;
parameter WEIGHT_0_2692 = 16'd2319;
parameter WEIGHT_0_2693 = 16'd4701;
parameter WEIGHT_0_2694 = 16'd-691;
parameter WEIGHT_0_2695 = 16'd-7959;
parameter WEIGHT_0_2696 = 16'd-15787;
parameter WEIGHT_0_2697 = 16'd10835;
parameter WEIGHT_0_2698 = 16'd-2975;
parameter WEIGHT_0_2699 = 16'd-3027;
parameter WEIGHT_0_2700 = 16'd6730;
parameter WEIGHT_0_2701 = 16'd-615;
parameter WEIGHT_0_2702 = 16'd1205;
parameter WEIGHT_0_2703 = 16'd4548;
parameter WEIGHT_0_2704 = 16'd-33;
parameter WEIGHT_0_2705 = 16'd-2304;
parameter WEIGHT_0_2706 = 16'd-15616;
parameter WEIGHT_0_2707 = 16'd5873;
parameter WEIGHT_0_2708 = 16'd1157;
parameter WEIGHT_0_2709 = 16'd-1975;
parameter WEIGHT_0_2710 = 16'd5222;
parameter WEIGHT_0_2711 = 16'd-6559;
parameter WEIGHT_0_2712 = 16'd-553;
parameter WEIGHT_0_2713 = 16'd4061;
parameter WEIGHT_0_2714 = 16'd-656;
parameter WEIGHT_0_2715 = 16'd-4532;
parameter WEIGHT_0_2716 = 16'd-11573;
parameter WEIGHT_0_2717 = 16'd7248;
parameter WEIGHT_0_2718 = 16'd2127;
parameter WEIGHT_0_2719 = 16'd-1408;
parameter WEIGHT_0_2720 = 16'd2310;
parameter WEIGHT_0_2721 = 16'd-7640;
parameter WEIGHT_0_2722 = 16'd454;
parameter WEIGHT_0_2723 = 16'd8054;
parameter WEIGHT_0_2724 = 16'd-1210;
parameter WEIGHT_0_2725 = 16'd912;
parameter WEIGHT_0_2726 = 16'd-7722;
parameter WEIGHT_0_2727 = 16'd3065;
parameter WEIGHT_0_2728 = 16'd3190;
parameter WEIGHT_0_2729 = 16'd-310;
parameter WEIGHT_0_2730 = 16'd3241;
parameter WEIGHT_0_2731 = 16'd-6515;
parameter WEIGHT_0_2732 = 16'd-763;
parameter WEIGHT_0_2733 = 16'd6241;
parameter WEIGHT_0_2734 = 16'd-2639;
parameter WEIGHT_0_2735 = 16'd6664;
parameter WEIGHT_0_2736 = 16'd-5063;
parameter WEIGHT_0_2737 = 16'd2416;
parameter WEIGHT_0_2738 = 16'd5440;
parameter WEIGHT_0_2739 = 16'd-3359;
parameter WEIGHT_0_2740 = 16'd3172;
parameter WEIGHT_0_2741 = 16'd-11698;
parameter WEIGHT_0_2742 = 16'd-10;
parameter WEIGHT_0_2743 = 16'd4179;
parameter WEIGHT_0_2744 = 16'd-3489;
parameter WEIGHT_0_2745 = 16'd9276;
parameter WEIGHT_0_2746 = 16'd-9795;
parameter WEIGHT_0_2747 = 16'd-338;
parameter WEIGHT_0_2748 = 16'd4850;
parameter WEIGHT_0_2749 = 16'd-6650;
parameter WEIGHT_0_2750 = 16'd3732;
parameter WEIGHT_0_2751 = 16'd-19293;
parameter WEIGHT_0_2752 = 16'd-8254;
parameter WEIGHT_0_2753 = 16'd-11760;
parameter WEIGHT_0_2754 = 16'd-3556;
parameter WEIGHT_0_2755 = 16'd14916;
parameter WEIGHT_0_2756 = 16'd-12005;
parameter WEIGHT_0_2757 = 16'd-5861;
parameter WEIGHT_0_2758 = 16'd2419;
parameter WEIGHT_0_2759 = 16'd-13456;
parameter WEIGHT_0_2760 = 16'd-1727;
parameter WEIGHT_0_2761 = 16'd-16234;
parameter WEIGHT_0_2762 = 16'd-26387;
parameter WEIGHT_0_2763 = 16'd-36087;
parameter WEIGHT_0_2764 = 16'd-14713;
parameter WEIGHT_0_2765 = 16'd24018;
parameter WEIGHT_0_2766 = 16'd-16044;
parameter WEIGHT_0_2767 = 16'd-12135;
parameter WEIGHT_0_2768 = 16'd-2224;
parameter WEIGHT_0_2769 = 16'd-17533;
parameter WEIGHT_0_2770 = 16'd-20336;
parameter WEIGHT_0_2771 = 16'd-17687;
parameter WEIGHT_0_2772 = 16'd-20045;
parameter WEIGHT_0_2773 = 16'd-14809;
parameter WEIGHT_0_2774 = 16'd-15030;
parameter WEIGHT_0_2775 = 16'd26982;
parameter WEIGHT_0_2776 = 16'd-25013;
parameter WEIGHT_0_2777 = 16'd-10960;
parameter WEIGHT_0_2778 = 16'd-4610;
parameter WEIGHT_0_2779 = 16'd-17372;
parameter WEIGHT_0_2780 = 16'd-18207;
parameter WEIGHT_0_2781 = 16'd-12142;
parameter WEIGHT_0_2782 = 16'd-5423;
parameter WEIGHT_0_2783 = 16'd-8368;
parameter WEIGHT_0_2784 = 16'd-12463;
parameter WEIGHT_0_2785 = 16'd10185;
parameter WEIGHT_0_2786 = 16'd-19128;
parameter WEIGHT_0_2787 = 16'd-7258;
parameter WEIGHT_0_2788 = 16'd2616;
parameter WEIGHT_0_2789 = 16'd-12630;
parameter WEIGHT_0_2790 = 16'd-6205;
parameter WEIGHT_0_2791 = 16'd-1457;
parameter WEIGHT_0_2792 = 16'd-4595;
parameter WEIGHT_0_2793 = 16'd-4249;
parameter WEIGHT_0_2794 = 16'd-4249;
parameter WEIGHT_0_2795 = 16'd4230;
parameter WEIGHT_0_2796 = 16'd-8640;
parameter WEIGHT_0_2797 = 16'd1460;
parameter WEIGHT_0_2798 = 16'd-2185;
parameter WEIGHT_0_2799 = 16'd-4317;
parameter WEIGHT_0_2800 = 16'd-3412;
parameter WEIGHT_0_2801 = 16'd-1396;
parameter WEIGHT_0_2802 = 16'd-3411;
parameter WEIGHT_0_2803 = 16'd-2780;
parameter WEIGHT_0_2804 = 16'd-3284;
parameter WEIGHT_0_2805 = 16'd-2557;
parameter WEIGHT_0_2806 = 16'd716;
parameter WEIGHT_0_2807 = 16'd5605;
parameter WEIGHT_0_2808 = 16'd-2347;
parameter WEIGHT_0_2809 = 16'd-2578;
parameter WEIGHT_0_2810 = 16'd313;
parameter WEIGHT_0_2811 = 16'd556;
parameter WEIGHT_0_2812 = 16'd-1063;
parameter WEIGHT_0_2813 = 16'd-2884;
parameter WEIGHT_0_2814 = 16'd-5724;
parameter WEIGHT_0_2815 = 16'd-2284;
parameter WEIGHT_0_2816 = 16'd-2614;
parameter WEIGHT_0_2817 = 16'd6326;
parameter WEIGHT_0_2818 = 16'd-1965;
parameter WEIGHT_0_2819 = 16'd-5938;
parameter WEIGHT_0_2820 = 16'd-1198;
parameter WEIGHT_0_2821 = 16'd-3609;
parameter WEIGHT_0_2822 = 16'd-154;
parameter WEIGHT_0_2823 = 16'd-422;
parameter WEIGHT_0_2824 = 16'd-7512;
parameter WEIGHT_0_2825 = 16'd-8677;
parameter WEIGHT_0_2826 = 16'd-4464;
parameter WEIGHT_0_2827 = 16'd10247;
parameter WEIGHT_0_2828 = 16'd-8965;
parameter WEIGHT_0_2829 = 16'd-12484;
parameter WEIGHT_0_2830 = 16'd-1181;
parameter WEIGHT_0_2831 = 16'd-2900;
parameter WEIGHT_0_2832 = 16'd4983;
parameter WEIGHT_0_2833 = 16'd6033;
parameter WEIGHT_0_2834 = 16'd-8413;
parameter WEIGHT_0_2835 = 16'd-11173;
parameter WEIGHT_0_2836 = 16'd-9264;
parameter WEIGHT_0_2837 = 16'd10561;
parameter WEIGHT_0_2838 = 16'd-5008;
parameter WEIGHT_0_2839 = 16'd-12055;
parameter WEIGHT_0_2840 = 16'd-4989;
parameter WEIGHT_0_2841 = 16'd-3705;
parameter WEIGHT_0_2842 = 16'd1956;
parameter WEIGHT_0_2843 = 16'd3607;
parameter WEIGHT_0_2844 = 16'd-8038;
parameter WEIGHT_0_2845 = 16'd-4359;
parameter WEIGHT_0_2846 = 16'd-8824;
parameter WEIGHT_0_2847 = 16'd9572;
parameter WEIGHT_0_2848 = 16'd1408;
parameter WEIGHT_0_2849 = 16'd-5776;
parameter WEIGHT_0_2850 = 16'd-1691;
parameter WEIGHT_0_2851 = 16'd-13088;
parameter WEIGHT_0_2852 = 16'd4785;
parameter WEIGHT_0_2853 = 16'd1075;
parameter WEIGHT_0_2854 = 16'd-8404;
parameter WEIGHT_0_2855 = 16'd-6696;
parameter WEIGHT_0_2856 = 16'd-8028;
parameter WEIGHT_0_2857 = 16'd3798;
parameter WEIGHT_0_2858 = 16'd1354;
parameter WEIGHT_0_2859 = 16'd-1435;
parameter WEIGHT_0_2860 = 16'd-4686;
parameter WEIGHT_0_2861 = 16'd-11017;
parameter WEIGHT_0_2862 = 16'd1989;
parameter WEIGHT_0_2863 = 16'd-2640;
parameter WEIGHT_0_2864 = 16'd-3881;
parameter WEIGHT_0_2865 = 16'd-621;
parameter WEIGHT_0_2866 = 16'd-2542;
parameter WEIGHT_0_2867 = 16'd-1424;
parameter WEIGHT_0_2868 = 16'd6325;
parameter WEIGHT_0_2869 = 16'd1763;
parameter WEIGHT_0_2870 = 16'd-2189;
parameter WEIGHT_0_2871 = 16'd-7732;
parameter WEIGHT_0_2872 = 16'd-6882;
parameter WEIGHT_0_2873 = 16'd-5187;
parameter WEIGHT_0_2874 = 16'd-3071;
parameter WEIGHT_0_2875 = 16'd4163;
parameter WEIGHT_0_2876 = 16'd-2483;
parameter WEIGHT_0_2877 = 16'd466;
parameter WEIGHT_0_2878 = 16'd3499;
parameter WEIGHT_0_2879 = 16'd-951;
parameter WEIGHT_0_2880 = 16'd-3746;
parameter WEIGHT_0_2881 = 16'd-6174;
parameter WEIGHT_0_2882 = 16'd-3671;
parameter WEIGHT_0_2883 = 16'd-11215;
parameter WEIGHT_0_2884 = 16'd-2785;
parameter WEIGHT_0_2885 = 16'd5961;
parameter WEIGHT_0_2886 = 16'd-1529;
parameter WEIGHT_0_2887 = 16'd-1421;
parameter WEIGHT_0_2888 = 16'd3626;
parameter WEIGHT_0_2889 = 16'd4059;
parameter WEIGHT_0_2890 = 16'd-2985;
parameter WEIGHT_0_2891 = 16'd-8455;
parameter WEIGHT_0_2892 = 16'd-5810;
parameter WEIGHT_0_2893 = 16'd-12866;
parameter WEIGHT_0_2894 = 16'd2852;
parameter WEIGHT_0_2895 = 16'd6970;
parameter WEIGHT_0_2896 = 16'd-1922;
parameter WEIGHT_0_2897 = 16'd422;
parameter WEIGHT_0_2898 = 16'd5792;
parameter WEIGHT_0_2899 = 16'd1459;
parameter WEIGHT_0_2900 = 16'd-1172;
parameter WEIGHT_0_2901 = 16'd-5909;
parameter WEIGHT_0_2902 = 16'd-2922;
parameter WEIGHT_0_2903 = 16'd-14516;
parameter WEIGHT_0_2904 = 16'd2348;
parameter WEIGHT_0_2905 = 16'd7151;
parameter WEIGHT_0_2906 = 16'd-4348;
parameter WEIGHT_0_2907 = 16'd79;
parameter WEIGHT_0_2908 = 16'd5461;
parameter WEIGHT_0_2909 = 16'd3449;
parameter WEIGHT_0_2910 = 16'd-2362;
parameter WEIGHT_0_2911 = 16'd345;
parameter WEIGHT_0_2912 = 16'd-6272;
parameter WEIGHT_0_2913 = 16'd-15066;
parameter WEIGHT_0_2914 = 16'd1357;
parameter WEIGHT_0_2915 = 16'd7446;
parameter WEIGHT_0_2916 = 16'd-3574;
parameter WEIGHT_0_2917 = 16'd861;
parameter WEIGHT_0_2918 = 16'd4938;
parameter WEIGHT_0_2919 = 16'd3744;
parameter WEIGHT_0_2920 = 16'd-791;
parameter WEIGHT_0_2921 = 16'd-3185;
parameter WEIGHT_0_2922 = 16'd-3780;
parameter WEIGHT_0_2923 = 16'd-10129;
parameter WEIGHT_0_2924 = 16'd1926;
parameter WEIGHT_0_2925 = 16'd6269;
parameter WEIGHT_0_2926 = 16'd-3345;
parameter WEIGHT_0_2927 = 16'd-688;
parameter WEIGHT_0_2928 = 16'd5072;
parameter WEIGHT_0_2929 = 16'd2379;
parameter WEIGHT_0_2930 = 16'd1797;
parameter WEIGHT_0_2931 = 16'd6167;
parameter WEIGHT_0_2932 = 16'd-7541;
parameter WEIGHT_0_2933 = 16'd-314;
parameter WEIGHT_0_2934 = 16'd-6442;
parameter WEIGHT_0_2935 = 16'd6720;
parameter WEIGHT_0_2936 = 16'd-2265;
parameter WEIGHT_0_2937 = 16'd6821;
parameter WEIGHT_0_2938 = 16'd474;
parameter WEIGHT_0_2939 = 16'd-2290;
parameter WEIGHT_0_2940 = 16'd-1267;
parameter WEIGHT_0_2941 = 16'd12749;
parameter WEIGHT_0_2942 = 16'd-3202;
parameter WEIGHT_0_2943 = 16'd2517;
parameter WEIGHT_0_2944 = 16'd-18872;
parameter WEIGHT_0_2945 = 16'd-1011;
parameter WEIGHT_0_2946 = 16'd-5052;
parameter WEIGHT_0_2947 = 16'd4665;
parameter WEIGHT_0_2948 = 16'd-3447;
parameter WEIGHT_0_2949 = 16'd-3326;
parameter WEIGHT_0_2950 = 16'd-3718;
parameter WEIGHT_0_2951 = 16'd12870;
parameter WEIGHT_0_2952 = 16'd-3925;
parameter WEIGHT_0_2953 = 16'd7014;
parameter WEIGHT_0_2954 = 16'd-8332;
parameter WEIGHT_0_2955 = 16'd-5160;
parameter WEIGHT_0_2956 = 16'd-9972;
parameter WEIGHT_0_2957 = 16'd12313;
parameter WEIGHT_0_2958 = 16'd-10031;
parameter WEIGHT_0_2959 = 16'd-5458;
parameter WEIGHT_0_2960 = 16'd-1676;
parameter WEIGHT_0_2961 = 16'd7450;
parameter WEIGHT_0_2962 = 16'd-127;
parameter WEIGHT_0_2963 = 16'd6553;
parameter WEIGHT_0_2964 = 16'd-2126;
parameter WEIGHT_0_2965 = 16'd-8705;
parameter WEIGHT_0_2966 = 16'd-14373;
parameter WEIGHT_0_2967 = 16'd11862;
parameter WEIGHT_0_2968 = 16'd-7083;
parameter WEIGHT_0_2969 = 16'd-2682;
parameter WEIGHT_0_2970 = 16'd4179;
parameter WEIGHT_0_2971 = 16'd-778;
parameter WEIGHT_0_2972 = 16'd-1232;
parameter WEIGHT_0_2973 = 16'd5196;
parameter WEIGHT_0_2974 = 16'd682;
parameter WEIGHT_0_2975 = 16'd-8338;
parameter WEIGHT_0_2976 = 16'd-13862;
parameter WEIGHT_0_2977 = 16'd9174;
parameter WEIGHT_0_2978 = 16'd-3425;
parameter WEIGHT_0_2979 = 16'd2379;
parameter WEIGHT_0_2980 = 16'd4895;
parameter WEIGHT_0_2981 = 16'd-5785;
parameter WEIGHT_0_2982 = 16'd-617;
parameter WEIGHT_0_2983 = 16'd5288;
parameter WEIGHT_0_2984 = 16'd-1255;
parameter WEIGHT_0_2985 = 16'd-10832;
parameter WEIGHT_0_2986 = 16'd-9208;
parameter WEIGHT_0_2987 = 16'd8863;
parameter WEIGHT_0_2988 = 16'd-998;
parameter WEIGHT_0_2989 = 16'd2244;
parameter WEIGHT_0_2990 = 16'd4294;
parameter WEIGHT_0_2991 = 16'd-6074;
parameter WEIGHT_0_2992 = 16'd-293;
parameter WEIGHT_0_2993 = 16'd2882;
parameter WEIGHT_0_2994 = 16'd-575;
parameter WEIGHT_0_2995 = 16'd-8349;
parameter WEIGHT_0_2996 = 16'd-9479;
parameter WEIGHT_0_2997 = 16'd6776;
parameter WEIGHT_0_2998 = 16'd2464;
parameter WEIGHT_0_2999 = 16'd207;
parameter WEIGHT_0_3000 = 16'd2856;
parameter WEIGHT_0_3001 = 16'd-7133;
parameter WEIGHT_0_3002 = 16'd655;
parameter WEIGHT_0_3003 = 16'd4082;
parameter WEIGHT_0_3004 = 16'd-952;
parameter WEIGHT_0_3005 = 16'd-6900;
parameter WEIGHT_0_3006 = 16'd-8712;
parameter WEIGHT_0_3007 = 16'd4880;
parameter WEIGHT_0_3008 = 16'd2489;
parameter WEIGHT_0_3009 = 16'd-931;
parameter WEIGHT_0_3010 = 16'd2225;
parameter WEIGHT_0_3011 = 16'd-11369;
parameter WEIGHT_0_3012 = 16'd-4437;
parameter WEIGHT_0_3013 = 16'd1926;
parameter WEIGHT_0_3014 = 16'd-2938;
parameter WEIGHT_0_3015 = 16'd-2353;
parameter WEIGHT_0_3016 = 16'd-5681;
parameter WEIGHT_0_3017 = 16'd6756;
parameter WEIGHT_0_3018 = 16'd3395;
parameter WEIGHT_0_3019 = 16'd-1717;
parameter WEIGHT_0_3020 = 16'd5644;
parameter WEIGHT_0_3021 = 16'd-15309;
parameter WEIGHT_0_3022 = 16'd-522;
parameter WEIGHT_0_3023 = 16'd-355;
parameter WEIGHT_0_3024 = 16'd-2282;
parameter WEIGHT_0_3025 = 16'd793;
parameter WEIGHT_0_3026 = 16'd-3870;
parameter WEIGHT_0_3027 = 16'd3979;
parameter WEIGHT_0_3028 = 16'd3362;
parameter WEIGHT_0_3029 = 16'd-1054;
parameter WEIGHT_0_3030 = 16'd9432;
parameter WEIGHT_0_3031 = 16'd-17632;
parameter WEIGHT_0_3032 = 16'd-3741;
parameter WEIGHT_0_3033 = 16'd-5879;
parameter WEIGHT_0_3034 = 16'd-11123;
parameter WEIGHT_0_3035 = 16'd11779;
parameter WEIGHT_0_3036 = 16'd-3798;
parameter WEIGHT_0_3037 = 16'd-3952;
parameter WEIGHT_0_3038 = 16'd3651;
parameter WEIGHT_0_3039 = 16'd-7434;
parameter WEIGHT_0_3040 = 16'd6191;
parameter WEIGHT_0_3041 = 16'd-25215;
parameter WEIGHT_0_3042 = 16'd-16210;
parameter WEIGHT_0_3043 = 16'd-25354;
parameter WEIGHT_0_3044 = 16'd-14363;
parameter WEIGHT_0_3045 = 16'd27123;
parameter WEIGHT_0_3046 = 16'd-9667;
parameter WEIGHT_0_3047 = 16'd-16218;
parameter WEIGHT_0_3048 = 16'd-6269;
parameter WEIGHT_0_3049 = 16'd-14163;
parameter WEIGHT_0_3050 = 16'd-15506;
parameter WEIGHT_0_3051 = 16'd-12073;
parameter WEIGHT_0_3052 = 16'd-7072;
parameter WEIGHT_0_3053 = 16'd-8215;
parameter WEIGHT_0_3054 = 16'd-13054;
parameter WEIGHT_0_3055 = 16'd28157;
parameter WEIGHT_0_3056 = 16'd-22882;
parameter WEIGHT_0_3057 = 16'd-10925;
parameter WEIGHT_0_3058 = 16'd-8945;
parameter WEIGHT_0_3059 = 16'd-14296;
parameter WEIGHT_0_3060 = 16'd-15086;
parameter WEIGHT_0_3061 = 16'd-7575;
parameter WEIGHT_0_3062 = 16'd489;
parameter WEIGHT_0_3063 = 16'd-4274;
parameter WEIGHT_0_3064 = 16'd-13638;
parameter WEIGHT_0_3065 = 16'd19513;
parameter WEIGHT_0_3066 = 16'd-16251;
parameter WEIGHT_0_3067 = 16'd-7343;
parameter WEIGHT_0_3068 = 16'd-3539;
parameter WEIGHT_0_3069 = 16'd-12165;
parameter WEIGHT_0_3070 = 16'd-3456;
parameter WEIGHT_0_3071 = 16'd-1589;
parameter WEIGHT_0_3072 = 16'd-3341;
parameter WEIGHT_0_3073 = 16'd-7245;
parameter WEIGHT_0_3074 = 16'd-3196;
parameter WEIGHT_0_3075 = 16'd5713;
parameter WEIGHT_0_3076 = 16'd-5401;
parameter WEIGHT_0_3077 = 16'd120;
parameter WEIGHT_0_3078 = 16'd2373;
parameter WEIGHT_0_3079 = 16'd-4629;
parameter WEIGHT_0_3080 = 16'd-3927;
parameter WEIGHT_0_3081 = 16'd691;
parameter WEIGHT_0_3082 = 16'd-871;
parameter WEIGHT_0_3083 = 16'd-6438;
parameter WEIGHT_0_3084 = 16'd-4275;
parameter WEIGHT_0_3085 = 16'd-4958;
parameter WEIGHT_0_3086 = 16'd1459;
parameter WEIGHT_0_3087 = 16'd1328;
parameter WEIGHT_0_3088 = 16'd-2953;
parameter WEIGHT_0_3089 = 16'd-1900;
parameter WEIGHT_0_3090 = 16'd2068;
parameter WEIGHT_0_3091 = 16'd3728;
parameter WEIGHT_0_3092 = 16'd-6437;
parameter WEIGHT_0_3093 = 16'd-6314;
parameter WEIGHT_0_3094 = 16'd-3407;
parameter WEIGHT_0_3095 = 16'd-9907;
parameter WEIGHT_0_3096 = 16'd-4835;
parameter WEIGHT_0_3097 = 16'd7376;
parameter WEIGHT_0_3098 = 16'd-5550;
parameter WEIGHT_0_3099 = 16'd-7354;
parameter WEIGHT_0_3100 = 16'd-680;
parameter WEIGHT_0_3101 = 16'd1147;
parameter WEIGHT_0_3102 = 16'd-3950;
parameter WEIGHT_0_3103 = 16'd558;
parameter WEIGHT_0_3104 = 16'd-9299;
parameter WEIGHT_0_3105 = 16'd-8949;
parameter WEIGHT_0_3106 = 16'd-418;
parameter WEIGHT_0_3107 = 16'd12300;
parameter WEIGHT_0_3108 = 16'd-11776;
parameter WEIGHT_0_3109 = 16'd-14257;
parameter WEIGHT_0_3110 = 16'd-2400;
parameter WEIGHT_0_3111 = 16'd-1434;
parameter WEIGHT_0_3112 = 16'd-1907;
parameter WEIGHT_0_3113 = 16'd9656;
parameter WEIGHT_0_3114 = 16'd-5033;
parameter WEIGHT_0_3115 = 16'd-11835;
parameter WEIGHT_0_3116 = 16'd-8187;
parameter WEIGHT_0_3117 = 16'd10003;
parameter WEIGHT_0_3118 = 16'd-7373;
parameter WEIGHT_0_3119 = 16'd-8847;
parameter WEIGHT_0_3120 = 16'd-7862;
parameter WEIGHT_0_3121 = 16'd-93;
parameter WEIGHT_0_3122 = 16'd-4488;
parameter WEIGHT_0_3123 = 16'd1167;
parameter WEIGHT_0_3124 = 16'd-5074;
parameter WEIGHT_0_3125 = 16'd-4396;
parameter WEIGHT_0_3126 = 16'd-3796;
parameter WEIGHT_0_3127 = 16'd9367;
parameter WEIGHT_0_3128 = 16'd244;
parameter WEIGHT_0_3129 = 16'd-3867;
parameter WEIGHT_0_3130 = 16'd-3520;
parameter WEIGHT_0_3131 = 16'd-8531;
parameter WEIGHT_0_3132 = 16'd-5451;
parameter WEIGHT_0_3133 = 16'd-4595;
parameter WEIGHT_0_3134 = 16'd-5267;
parameter WEIGHT_0_3135 = 16'd-1517;
parameter WEIGHT_0_3136 = 16'd-1635;
parameter WEIGHT_0_3137 = 16'd4246;
parameter WEIGHT_0_3138 = 16'd2076;
parameter WEIGHT_0_3139 = 16'd6949;
parameter WEIGHT_0_3140 = 16'd-2543;
parameter WEIGHT_0_3141 = 16'd-12023;
parameter WEIGHT_0_3142 = 16'd-5533;
parameter WEIGHT_0_3143 = 16'd-6852;
parameter WEIGHT_0_3144 = 16'd-532;
parameter WEIGHT_0_3145 = 16'd4790;
parameter WEIGHT_0_3146 = 16'd-1314;
parameter WEIGHT_0_3147 = 16'd49;
parameter WEIGHT_0_3148 = 16'd3778;
parameter WEIGHT_0_3149 = 16'd6852;
parameter WEIGHT_0_3150 = 16'd387;
parameter WEIGHT_0_3151 = 16'd-5082;
parameter WEIGHT_0_3152 = 16'd-11439;
parameter WEIGHT_0_3153 = 16'd-11857;
parameter WEIGHT_0_3154 = 16'd304;
parameter WEIGHT_0_3155 = 16'd3738;
parameter WEIGHT_0_3156 = 16'd4383;
parameter WEIGHT_0_3157 = 16'd832;
parameter WEIGHT_0_3158 = 16'd4916;
parameter WEIGHT_0_3159 = 16'd3525;
parameter WEIGHT_0_3160 = 16'd-2022;
parameter WEIGHT_0_3161 = 16'd-5190;
parameter WEIGHT_0_3162 = 16'd-11458;
parameter WEIGHT_0_3163 = 16'd-12540;
parameter WEIGHT_0_3164 = 16'd493;
parameter WEIGHT_0_3165 = 16'd4914;
parameter WEIGHT_0_3166 = 16'd-1523;
parameter WEIGHT_0_3167 = 16'd248;
parameter WEIGHT_0_3168 = 16'd8942;
parameter WEIGHT_0_3169 = 16'd4339;
parameter WEIGHT_0_3170 = 16'd-3856;
parameter WEIGHT_0_3171 = 16'd-6876;
parameter WEIGHT_0_3172 = 16'd-10919;
parameter WEIGHT_0_3173 = 16'd-14451;
parameter WEIGHT_0_3174 = 16'd6145;
parameter WEIGHT_0_3175 = 16'd2041;
parameter WEIGHT_0_3176 = 16'd3199;
parameter WEIGHT_0_3177 = 16'd646;
parameter WEIGHT_0_3178 = 16'd5627;
parameter WEIGHT_0_3179 = 16'd3360;
parameter WEIGHT_0_3180 = 16'd-1366;
parameter WEIGHT_0_3181 = 16'd-4144;
parameter WEIGHT_0_3182 = 16'd-16176;
parameter WEIGHT_0_3183 = 16'd-9712;
parameter WEIGHT_0_3184 = 16'd5186;
parameter WEIGHT_0_3185 = 16'd2834;
parameter WEIGHT_0_3186 = 16'd1522;
parameter WEIGHT_0_3187 = 16'd3186;
parameter WEIGHT_0_3188 = 16'd3282;
parameter WEIGHT_0_3189 = 16'd5609;
parameter WEIGHT_0_3190 = 16'd732;
parameter WEIGHT_0_3191 = 16'd-6525;
parameter WEIGHT_0_3192 = 16'd-15468;
parameter WEIGHT_0_3193 = 16'd-6915;
parameter WEIGHT_0_3194 = 16'd9021;
parameter WEIGHT_0_3195 = 16'd6577;
parameter WEIGHT_0_3196 = 16'd893;
parameter WEIGHT_0_3197 = 16'd1417;
parameter WEIGHT_0_3198 = 16'd1831;
parameter WEIGHT_0_3199 = 16'd2444;
parameter WEIGHT_0_3200 = 16'd-193;
parameter WEIGHT_0_3201 = 16'd-5733;
parameter WEIGHT_0_3202 = 16'd-21278;
parameter WEIGHT_0_3203 = 16'd-5586;
parameter WEIGHT_0_3204 = 16'd5294;
parameter WEIGHT_0_3205 = 16'd9163;
parameter WEIGHT_0_3206 = 16'd-638;
parameter WEIGHT_0_3207 = 16'd-3412;
parameter WEIGHT_0_3208 = 16'd2812;
parameter WEIGHT_0_3209 = 16'd-2987;
parameter WEIGHT_0_3210 = 16'd-6202;
parameter WEIGHT_0_3211 = 16'd5783;
parameter WEIGHT_0_3212 = 16'd-22335;
parameter WEIGHT_0_3213 = 16'd2943;
parameter WEIGHT_0_3214 = 16'd-10826;
parameter WEIGHT_0_3215 = 16'd10545;
parameter WEIGHT_0_3216 = 16'd2132;
parameter WEIGHT_0_3217 = 16'd-851;
parameter WEIGHT_0_3218 = 16'd5575;
parameter WEIGHT_0_3219 = 16'd-3567;
parameter WEIGHT_0_3220 = 16'd-12604;
parameter WEIGHT_0_3221 = 16'd18370;
parameter WEIGHT_0_3222 = 16'd-17461;
parameter WEIGHT_0_3223 = 16'd4556;
parameter WEIGHT_0_3224 = 16'd-20034;
parameter WEIGHT_0_3225 = 16'd1234;
parameter WEIGHT_0_3226 = 16'd-5597;
parameter WEIGHT_0_3227 = 16'd4613;
parameter WEIGHT_0_3228 = 16'd6426;
parameter WEIGHT_0_3229 = 16'd-5116;
parameter WEIGHT_0_3230 = 16'd-15855;
parameter WEIGHT_0_3231 = 16'd18083;
parameter WEIGHT_0_3232 = 16'd-9745;
parameter WEIGHT_0_3233 = 16'd5579;
parameter WEIGHT_0_3234 = 16'd-2020;
parameter WEIGHT_0_3235 = 16'd-3183;
parameter WEIGHT_0_3236 = 16'd-15949;
parameter WEIGHT_0_3237 = 16'd11731;
parameter WEIGHT_0_3238 = 16'd-2772;
parameter WEIGHT_0_3239 = 16'd2929;
parameter WEIGHT_0_3240 = 16'd-16362;
parameter WEIGHT_0_3241 = 16'd6895;
parameter WEIGHT_0_3242 = 16'd-4670;
parameter WEIGHT_0_3243 = 16'd549;
parameter WEIGHT_0_3244 = 16'd7802;
parameter WEIGHT_0_3245 = 16'd-5415;
parameter WEIGHT_0_3246 = 16'd-9463;
parameter WEIGHT_0_3247 = 16'd10798;
parameter WEIGHT_0_3248 = 16'd-7476;
parameter WEIGHT_0_3249 = 16'd2153;
parameter WEIGHT_0_3250 = 16'd-3788;
parameter WEIGHT_0_3251 = 16'd-3823;
parameter WEIGHT_0_3252 = 16'd-3204;
parameter WEIGHT_0_3253 = 16'd2555;
parameter WEIGHT_0_3254 = 16'd2383;
parameter WEIGHT_0_3255 = 16'd-6245;
parameter WEIGHT_0_3256 = 16'd-9589;
parameter WEIGHT_0_3257 = 16'd12098;
parameter WEIGHT_0_3258 = 16'd-2716;
parameter WEIGHT_0_3259 = 16'd5211;
parameter WEIGHT_0_3260 = 16'd-1377;
parameter WEIGHT_0_3261 = 16'd-1188;
parameter WEIGHT_0_3262 = 16'd-2183;
parameter WEIGHT_0_3263 = 16'd2581;
parameter WEIGHT_0_3264 = 16'd1554;
parameter WEIGHT_0_3265 = 16'd-9082;
parameter WEIGHT_0_3266 = 16'd-8331;
parameter WEIGHT_0_3267 = 16'd9033;
parameter WEIGHT_0_3268 = 16'd-1668;
parameter WEIGHT_0_3269 = 16'd4967;
parameter WEIGHT_0_3270 = 16'd5084;
parameter WEIGHT_0_3271 = 16'd-2588;
parameter WEIGHT_0_3272 = 16'd2069;
parameter WEIGHT_0_3273 = 16'd5639;
parameter WEIGHT_0_3274 = 16'd-298;
parameter WEIGHT_0_3275 = 16'd-9625;
parameter WEIGHT_0_3276 = 16'd-3445;
parameter WEIGHT_0_3277 = 16'd3228;
parameter WEIGHT_0_3278 = 16'd486;
parameter WEIGHT_0_3279 = 16'd7219;
parameter WEIGHT_0_3280 = 16'd3794;
parameter WEIGHT_0_3281 = 16'd-7236;
parameter WEIGHT_0_3282 = 16'd403;
parameter WEIGHT_0_3283 = 16'd3473;
parameter WEIGHT_0_3284 = 16'd-3754;
parameter WEIGHT_0_3285 = 16'd-13765;
parameter WEIGHT_0_3286 = 16'd-2794;
parameter WEIGHT_0_3287 = 16'd5158;
parameter WEIGHT_0_3288 = 16'd2689;
parameter WEIGHT_0_3289 = 16'd9727;
parameter WEIGHT_0_3290 = 16'd7236;
parameter WEIGHT_0_3291 = 16'd-7881;
parameter WEIGHT_0_3292 = 16'd-4590;
parameter WEIGHT_0_3293 = 16'd-4209;
parameter WEIGHT_0_3294 = 16'd-2725;
parameter WEIGHT_0_3295 = 16'd-14368;
parameter WEIGHT_0_3296 = 16'd2972;
parameter WEIGHT_0_3297 = 16'd1937;
parameter WEIGHT_0_3298 = 16'd3734;
parameter WEIGHT_0_3299 = 16'd9027;
parameter WEIGHT_0_3300 = 16'd7562;
parameter WEIGHT_0_3301 = 16'd-10159;
parameter WEIGHT_0_3302 = 16'd-2371;
parameter WEIGHT_0_3303 = 16'd-2806;
parameter WEIGHT_0_3304 = 16'd-5281;
parameter WEIGHT_0_3305 = 16'd-12811;
parameter WEIGHT_0_3306 = 16'd1564;
parameter WEIGHT_0_3307 = 16'd1480;
parameter WEIGHT_0_3308 = 16'd9037;
parameter WEIGHT_0_3309 = 16'd3590;
parameter WEIGHT_0_3310 = 16'd6969;
parameter WEIGHT_0_3311 = 16'd-9956;
parameter WEIGHT_0_3312 = 16'd-8118;
parameter WEIGHT_0_3313 = 16'd-9795;
parameter WEIGHT_0_3314 = 16'd-13548;
parameter WEIGHT_0_3315 = 16'd-4131;
parameter WEIGHT_0_3316 = 16'd4806;
parameter WEIGHT_0_3317 = 16'd-5261;
parameter WEIGHT_0_3318 = 16'd7110;
parameter WEIGHT_0_3319 = 16'd-1766;
parameter WEIGHT_0_3320 = 16'd4731;
parameter WEIGHT_0_3321 = 16'd-13729;
parameter WEIGHT_0_3322 = 16'd-6825;
parameter WEIGHT_0_3323 = 16'd-19203;
parameter WEIGHT_0_3324 = 16'd-16947;
parameter WEIGHT_0_3325 = 16'd10492;
parameter WEIGHT_0_3326 = 16'd1709;
parameter WEIGHT_0_3327 = 16'd-15695;
parameter WEIGHT_0_3328 = 16'd5662;
parameter WEIGHT_0_3329 = 16'd-12908;
parameter WEIGHT_0_3330 = 16'd-11851;
parameter WEIGHT_0_3331 = 16'd-2286;
parameter WEIGHT_0_3332 = 16'd1375;
parameter WEIGHT_0_3333 = 16'd-5669;
parameter WEIGHT_0_3334 = 16'd-14881;
parameter WEIGHT_0_3335 = 16'd21620;
parameter WEIGHT_0_3336 = 16'd-10278;
parameter WEIGHT_0_3337 = 16'd-15076;
parameter WEIGHT_0_3338 = 16'd-238;
parameter WEIGHT_0_3339 = 16'd-14997;
parameter WEIGHT_0_3340 = 16'd-15425;
parameter WEIGHT_0_3341 = 16'd-2313;
parameter WEIGHT_0_3342 = 16'd936;
parameter WEIGHT_0_3343 = 16'd-5428;
parameter WEIGHT_0_3344 = 16'd-7998;
parameter WEIGHT_0_3345 = 16'd13547;
parameter WEIGHT_0_3346 = 16'd-16622;
parameter WEIGHT_0_3347 = 16'd-4623;
parameter WEIGHT_0_3348 = 16'd2202;
parameter WEIGHT_0_3349 = 16'd-10249;
parameter WEIGHT_0_3350 = 16'd-4746;
parameter WEIGHT_0_3351 = 16'd-668;
parameter WEIGHT_0_3352 = 16'd-4744;
parameter WEIGHT_0_3353 = 16'd-2762;
parameter WEIGHT_0_3354 = 16'd-3481;
parameter WEIGHT_0_3355 = 16'd2305;
parameter WEIGHT_0_3356 = 16'd-793;
parameter WEIGHT_0_3357 = 16'd-2232;
parameter WEIGHT_0_3358 = 16'd3094;
parameter WEIGHT_0_3359 = 16'd-5511;
parameter WEIGHT_0_3360 = 16'd972;
parameter WEIGHT_0_3361 = 16'd1392;
parameter WEIGHT_0_3362 = 16'd-3799;
parameter WEIGHT_0_3363 = 16'd-1350;
parameter WEIGHT_0_3364 = 16'd-1356;
parameter WEIGHT_0_3365 = 16'd-3052;
parameter WEIGHT_0_3366 = 16'd-2234;
parameter WEIGHT_0_3367 = 16'd-74;
parameter WEIGHT_0_3368 = 16'd-1271;
parameter WEIGHT_0_3369 = 16'd-3323;
parameter WEIGHT_0_3370 = 16'd-1723;
parameter WEIGHT_0_3371 = 16'd-3048;
parameter WEIGHT_0_3372 = 16'd-3080;
parameter WEIGHT_0_3373 = 16'd-7642;
parameter WEIGHT_0_3374 = 16'd-3908;
parameter WEIGHT_0_3375 = 16'd-4496;
parameter WEIGHT_0_3376 = 16'd-2235;
parameter WEIGHT_0_3377 = 16'd10924;
parameter WEIGHT_0_3378 = 16'd-8167;
parameter WEIGHT_0_3379 = 16'd-8659;
parameter WEIGHT_0_3380 = 16'd-4962;
parameter WEIGHT_0_3381 = 16'd-1044;
parameter WEIGHT_0_3382 = 16'd-1621;
parameter WEIGHT_0_3383 = 16'd-4488;
parameter WEIGHT_0_3384 = 16'd-10013;
parameter WEIGHT_0_3385 = 16'd-6371;
parameter WEIGHT_0_3386 = 16'd-674;
parameter WEIGHT_0_3387 = 16'd11880;
parameter WEIGHT_0_3388 = 16'd-11366;
parameter WEIGHT_0_3389 = 16'd-11996;
parameter WEIGHT_0_3390 = 16'd-5590;
parameter WEIGHT_0_3391 = 16'd-2725;
parameter WEIGHT_0_3392 = 16'd-5326;
parameter WEIGHT_0_3393 = 16'd-389;
parameter WEIGHT_0_3394 = 16'd-7774;
parameter WEIGHT_0_3395 = 16'd-4243;
parameter WEIGHT_0_3396 = 16'd-10616;
parameter WEIGHT_0_3397 = 16'd14302;
parameter WEIGHT_0_3398 = 16'd-2192;
parameter WEIGHT_0_3399 = 16'd-4238;
parameter WEIGHT_0_3400 = 16'd-4803;
parameter WEIGHT_0_3401 = 16'd-456;
parameter WEIGHT_0_3402 = 16'd-9696;
parameter WEIGHT_0_3403 = 16'd-3307;
parameter WEIGHT_0_3404 = 16'd-5014;
parameter WEIGHT_0_3405 = 16'd431;
parameter WEIGHT_0_3406 = 16'd-3760;
parameter WEIGHT_0_3407 = 16'd7901;
parameter WEIGHT_0_3408 = 16'd2958;
parameter WEIGHT_0_3409 = 16'd5450;
parameter WEIGHT_0_3410 = 16'd413;
parameter WEIGHT_0_3411 = 16'd-4510;
parameter WEIGHT_0_3412 = 16'd-11978;
parameter WEIGHT_0_3413 = 16'd-7751;
parameter WEIGHT_0_3414 = 16'd-767;
parameter WEIGHT_0_3415 = 16'd4240;
parameter WEIGHT_0_3416 = 16'd-2787;
parameter WEIGHT_0_3417 = 16'd2270;
parameter WEIGHT_0_3418 = 16'd4570;
parameter WEIGHT_0_3419 = 16'd8761;
parameter WEIGHT_0_3420 = 16'd902;
parameter WEIGHT_0_3421 = 16'd-3699;
parameter WEIGHT_0_3422 = 16'd-22620;
parameter WEIGHT_0_3423 = 16'd-11427;
parameter WEIGHT_0_3424 = 16'd664;
parameter WEIGHT_0_3425 = 16'd6264;
parameter WEIGHT_0_3426 = 16'd989;
parameter WEIGHT_0_3427 = 16'd429;
parameter WEIGHT_0_3428 = 16'd5167;
parameter WEIGHT_0_3429 = 16'd6955;
parameter WEIGHT_0_3430 = 16'd19;
parameter WEIGHT_0_3431 = 16'd-4665;
parameter WEIGHT_0_3432 = 16'd-20798;
parameter WEIGHT_0_3433 = 16'd-12493;
parameter WEIGHT_0_3434 = 16'd6742;
parameter WEIGHT_0_3435 = 16'd1974;
parameter WEIGHT_0_3436 = 16'd2489;
parameter WEIGHT_0_3437 = 16'd2419;
parameter WEIGHT_0_3438 = 16'd3821;
parameter WEIGHT_0_3439 = 16'd6747;
parameter WEIGHT_0_3440 = 16'd212;
parameter WEIGHT_0_3441 = 16'd-3730;
parameter WEIGHT_0_3442 = 16'd-16965;
parameter WEIGHT_0_3443 = 16'd-10488;
parameter WEIGHT_0_3444 = 16'd7406;
parameter WEIGHT_0_3445 = 16'd3009;
parameter WEIGHT_0_3446 = 16'd2956;
parameter WEIGHT_0_3447 = 16'd3231;
parameter WEIGHT_0_3448 = 16'd2656;
parameter WEIGHT_0_3449 = 16'd5076;
parameter WEIGHT_0_3450 = 16'd-3523;
parameter WEIGHT_0_3451 = 16'd-5240;
parameter WEIGHT_0_3452 = 16'd-17369;
parameter WEIGHT_0_3453 = 16'd-5988;
parameter WEIGHT_0_3454 = 16'd7189;
parameter WEIGHT_0_3455 = 16'd-964;
parameter WEIGHT_0_3456 = 16'd1507;
parameter WEIGHT_0_3457 = 16'd-1767;
parameter WEIGHT_0_3458 = 16'd3551;
parameter WEIGHT_0_3459 = 16'd6285;
parameter WEIGHT_0_3460 = 16'd-3383;
parameter WEIGHT_0_3461 = 16'd-10151;
parameter WEIGHT_0_3462 = 16'd-16856;
parameter WEIGHT_0_3463 = 16'd-4086;
parameter WEIGHT_0_3464 = 16'd8933;
parameter WEIGHT_0_3465 = 16'd5557;
parameter WEIGHT_0_3466 = 16'd687;
parameter WEIGHT_0_3467 = 16'd-1716;
parameter WEIGHT_0_3468 = 16'd-885;
parameter WEIGHT_0_3469 = 16'd6260;
parameter WEIGHT_0_3470 = 16'd-2515;
parameter WEIGHT_0_3471 = 16'd-11197;
parameter WEIGHT_0_3472 = 16'd-18017;
parameter WEIGHT_0_3473 = 16'd-3720;
parameter WEIGHT_0_3474 = 16'd14245;
parameter WEIGHT_0_3475 = 16'd8478;
parameter WEIGHT_0_3476 = 16'd4981;
parameter WEIGHT_0_3477 = 16'd-6944;
parameter WEIGHT_0_3478 = 16'd-2245;
parameter WEIGHT_0_3479 = 16'd1880;
parameter WEIGHT_0_3480 = 16'd-2064;
parameter WEIGHT_0_3481 = 16'd-7669;
parameter WEIGHT_0_3482 = 16'd-17281;
parameter WEIGHT_0_3483 = 16'd-1528;
parameter WEIGHT_0_3484 = 16'd9553;
parameter WEIGHT_0_3485 = 16'd7124;
parameter WEIGHT_0_3486 = 16'd1982;
parameter WEIGHT_0_3487 = 16'd-14361;
parameter WEIGHT_0_3488 = 16'd3218;
parameter WEIGHT_0_3489 = 16'd-7058;
parameter WEIGHT_0_3490 = 16'd-5133;
parameter WEIGHT_0_3491 = 16'd6679;
parameter WEIGHT_0_3492 = 16'd-15767;
parameter WEIGHT_0_3493 = 16'd3009;
parameter WEIGHT_0_3494 = 16'd-5055;
parameter WEIGHT_0_3495 = 16'd6347;
parameter WEIGHT_0_3496 = 16'd379;
parameter WEIGHT_0_3497 = 16'd-14422;
parameter WEIGHT_0_3498 = 16'd7231;
parameter WEIGHT_0_3499 = 16'd-345;
parameter WEIGHT_0_3500 = 16'd-17639;
parameter WEIGHT_0_3501 = 16'd15784;
parameter WEIGHT_0_3502 = 16'd-12448;
parameter WEIGHT_0_3503 = 16'd5493;
parameter WEIGHT_0_3504 = 16'd-11463;
parameter WEIGHT_0_3505 = 16'd-474;
parameter WEIGHT_0_3506 = 16'd-9400;
parameter WEIGHT_0_3507 = 16'd-9937;
parameter WEIGHT_0_3508 = 16'd2312;
parameter WEIGHT_0_3509 = 16'd4084;
parameter WEIGHT_0_3510 = 16'd-20596;
parameter WEIGHT_0_3511 = 16'd15605;
parameter WEIGHT_0_3512 = 16'd-9800;
parameter WEIGHT_0_3513 = 16'd2072;
parameter WEIGHT_0_3514 = 16'd2777;
parameter WEIGHT_0_3515 = 16'd-6848;
parameter WEIGHT_0_3516 = 16'd-9965;
parameter WEIGHT_0_3517 = 16'd3842;
parameter WEIGHT_0_3518 = 16'd1903;
parameter WEIGHT_0_3519 = 16'd5124;
parameter WEIGHT_0_3520 = 16'd-16651;
parameter WEIGHT_0_3521 = 16'd5148;
parameter WEIGHT_0_3522 = 16'd-11242;
parameter WEIGHT_0_3523 = 16'd2195;
parameter WEIGHT_0_3524 = 16'd9132;
parameter WEIGHT_0_3525 = 16'd-11198;
parameter WEIGHT_0_3526 = 16'd-1649;
parameter WEIGHT_0_3527 = 16'd7197;
parameter WEIGHT_0_3528 = 16'd-1565;
parameter WEIGHT_0_3529 = 16'd6568;
parameter WEIGHT_0_3530 = 16'd-5830;
parameter WEIGHT_0_3531 = 16'd-1927;
parameter WEIGHT_0_3532 = 16'd-7106;
parameter WEIGHT_0_3533 = 16'd2336;
parameter WEIGHT_0_3534 = 16'd5226;
parameter WEIGHT_0_3535 = 16'd-10078;
parameter WEIGHT_0_3536 = 16'd-3126;
parameter WEIGHT_0_3537 = 16'd7699;
parameter WEIGHT_0_3538 = 16'd-3161;
parameter WEIGHT_0_3539 = 16'd11619;
parameter WEIGHT_0_3540 = 16'd-4729;
parameter WEIGHT_0_3541 = 16'd-4372;
parameter WEIGHT_0_3542 = 16'd-2825;
parameter WEIGHT_0_3543 = 16'd3307;
parameter WEIGHT_0_3544 = 16'd405;
parameter WEIGHT_0_3545 = 16'd-7259;
parameter WEIGHT_0_3546 = 16'd-4510;
parameter WEIGHT_0_3547 = 16'd6495;
parameter WEIGHT_0_3548 = 16'd402;
parameter WEIGHT_0_3549 = 16'd8661;
parameter WEIGHT_0_3550 = 16'd284;
parameter WEIGHT_0_3551 = 16'd-6841;
parameter WEIGHT_0_3552 = 16'd-2326;
parameter WEIGHT_0_3553 = 16'd-1180;
parameter WEIGHT_0_3554 = 16'd-287;
parameter WEIGHT_0_3555 = 16'd-9083;
parameter WEIGHT_0_3556 = 16'd-6524;
parameter WEIGHT_0_3557 = 16'd-503;
parameter WEIGHT_0_3558 = 16'd1940;
parameter WEIGHT_0_3559 = 16'd7565;
parameter WEIGHT_0_3560 = 16'd-462;
parameter WEIGHT_0_3561 = 16'd-4473;
parameter WEIGHT_0_3562 = 16'd-308;
parameter WEIGHT_0_3563 = 16'd-6164;
parameter WEIGHT_0_3564 = 16'd681;
parameter WEIGHT_0_3565 = 16'd-13264;
parameter WEIGHT_0_3566 = 16'd-2391;
parameter WEIGHT_0_3567 = 16'd-612;
parameter WEIGHT_0_3568 = 16'd4081;
parameter WEIGHT_0_3569 = 16'd7384;
parameter WEIGHT_0_3570 = 16'd1027;
parameter WEIGHT_0_3571 = 16'd-6310;
parameter WEIGHT_0_3572 = 16'd-1371;
parameter WEIGHT_0_3573 = 16'd-12884;
parameter WEIGHT_0_3574 = 16'd2528;
parameter WEIGHT_0_3575 = 16'd-21561;
parameter WEIGHT_0_3576 = 16'd4649;
parameter WEIGHT_0_3577 = 16'd-753;
parameter WEIGHT_0_3578 = 16'd5266;
parameter WEIGHT_0_3579 = 16'd8038;
parameter WEIGHT_0_3580 = 16'd6239;
parameter WEIGHT_0_3581 = 16'd-6931;
parameter WEIGHT_0_3582 = 16'd-5854;
parameter WEIGHT_0_3583 = 16'd-12803;
parameter WEIGHT_0_3584 = 16'd-869;
parameter WEIGHT_0_3585 = 16'd-25174;
parameter WEIGHT_0_3586 = 16'd8937;
parameter WEIGHT_0_3587 = 16'd-3362;
parameter WEIGHT_0_3588 = 16'd8313;
parameter WEIGHT_0_3589 = 16'd5169;
parameter WEIGHT_0_3590 = 16'd10934;
parameter WEIGHT_0_3591 = 16'd-5230;
parameter WEIGHT_0_3592 = 16'd-7148;
parameter WEIGHT_0_3593 = 16'd-12451;
parameter WEIGHT_0_3594 = 16'd-8787;
parameter WEIGHT_0_3595 = 16'd-24204;
parameter WEIGHT_0_3596 = 16'd12601;
parameter WEIGHT_0_3597 = 16'd-3752;
parameter WEIGHT_0_3598 = 16'd11589;
parameter WEIGHT_0_3599 = 16'd3990;
parameter WEIGHT_0_3600 = 16'd9287;
parameter WEIGHT_0_3601 = 16'd-11791;
parameter WEIGHT_0_3602 = 16'd-1609;
parameter WEIGHT_0_3603 = 16'd-16745;
parameter WEIGHT_0_3604 = 16'd-4912;
parameter WEIGHT_0_3605 = 16'd-18743;
parameter WEIGHT_0_3606 = 16'd5520;
parameter WEIGHT_0_3607 = 16'd-7925;
parameter WEIGHT_0_3608 = 16'd7582;
parameter WEIGHT_0_3609 = 16'd-15206;
parameter WEIGHT_0_3610 = 16'd-189;
parameter WEIGHT_0_3611 = 16'd-6538;
parameter WEIGHT_0_3612 = 16'd8913;
parameter WEIGHT_0_3613 = 16'd188;
parameter WEIGHT_0_3614 = 16'd-4024;
parameter WEIGHT_0_3615 = 16'd1003;
parameter WEIGHT_0_3616 = 16'd-5917;
parameter WEIGHT_0_3617 = 16'd-529;
parameter WEIGHT_0_3618 = 16'd1544;
parameter WEIGHT_0_3619 = 16'd-18372;
parameter WEIGHT_0_3620 = 16'd-9472;
parameter WEIGHT_0_3621 = 16'd-6826;
parameter WEIGHT_0_3622 = 16'd9917;
parameter WEIGHT_0_3623 = 16'd-4390;
parameter WEIGHT_0_3624 = 16'd-4527;
parameter WEIGHT_0_3625 = 16'd2059;
parameter WEIGHT_0_3626 = 16'd-12814;
parameter WEIGHT_0_3627 = 16'd-91;
parameter WEIGHT_0_3628 = 16'd953;
parameter WEIGHT_0_3629 = 16'd-14662;
parameter WEIGHT_0_3630 = 16'd-3266;
parameter WEIGHT_0_3631 = 16'd691;
parameter WEIGHT_0_3632 = 16'd3055;
parameter WEIGHT_0_3633 = 16'd-2011;
parameter WEIGHT_0_3634 = 16'd-8180;
parameter WEIGHT_0_3635 = 16'd-4113;
parameter WEIGHT_0_3636 = 16'd-4303;
parameter WEIGHT_0_3637 = 16'd2505;
parameter WEIGHT_0_3638 = 16'd-2250;
parameter WEIGHT_0_3639 = 16'd-3432;
parameter WEIGHT_0_3640 = 16'd98;
parameter WEIGHT_0_3641 = 16'd587;
parameter WEIGHT_0_3642 = 16'd-1329;
parameter WEIGHT_0_3643 = 16'd-3175;
parameter WEIGHT_0_3644 = 16'd1152;
parameter WEIGHT_0_3645 = 16'd-1271;
parameter WEIGHT_0_3646 = 16'd180;
parameter WEIGHT_0_3647 = 16'd-2338;
parameter WEIGHT_0_3648 = 16'd501;
parameter WEIGHT_0_3649 = 16'd-519;
parameter WEIGHT_0_3650 = 16'd2951;
parameter WEIGHT_0_3651 = 16'd50;
parameter WEIGHT_0_3652 = 16'd-64;
parameter WEIGHT_0_3653 = 16'd-5589;
parameter WEIGHT_0_3654 = 16'd-1426;
parameter WEIGHT_0_3655 = 16'd-2858;
parameter WEIGHT_0_3656 = 16'd-400;
parameter WEIGHT_0_3657 = 16'd6444;
parameter WEIGHT_0_3658 = 16'd-5250;
parameter WEIGHT_0_3659 = 16'd-2922;
parameter WEIGHT_0_3660 = 16'd1080;
parameter WEIGHT_0_3661 = 16'd-827;
parameter WEIGHT_0_3662 = 16'd506;
parameter WEIGHT_0_3663 = 16'd-9282;
parameter WEIGHT_0_3664 = 16'd-4659;
parameter WEIGHT_0_3665 = 16'd-8221;
parameter WEIGHT_0_3666 = 16'd-3420;
parameter WEIGHT_0_3667 = 16'd10957;
parameter WEIGHT_0_3668 = 16'd-5707;
parameter WEIGHT_0_3669 = 16'd-8592;
parameter WEIGHT_0_3670 = 16'd-1683;
parameter WEIGHT_0_3671 = 16'd784;
parameter WEIGHT_0_3672 = 16'd-6837;
parameter WEIGHT_0_3673 = 16'd-395;
parameter WEIGHT_0_3674 = 16'd-8987;
parameter WEIGHT_0_3675 = 16'd-2209;
parameter WEIGHT_0_3676 = 16'd-10860;
parameter WEIGHT_0_3677 = 16'd12100;
parameter WEIGHT_0_3678 = 16'd-4597;
parameter WEIGHT_0_3679 = 16'd-2023;
parameter WEIGHT_0_3680 = 16'd-4240;
parameter WEIGHT_0_3681 = 16'd-1267;
parameter WEIGHT_0_3682 = 16'd-15248;
parameter WEIGHT_0_3683 = 16'd-7877;
parameter WEIGHT_0_3684 = 16'd-4355;
parameter WEIGHT_0_3685 = 16'd2581;
parameter WEIGHT_0_3686 = 16'd-5289;
parameter WEIGHT_0_3687 = 16'd6221;
parameter WEIGHT_0_3688 = 16'd-839;
parameter WEIGHT_0_3689 = 16'd7608;
parameter WEIGHT_0_3690 = 16'd2040;
parameter WEIGHT_0_3691 = 16'd-5998;
parameter WEIGHT_0_3692 = 16'd-21859;
parameter WEIGHT_0_3693 = 16'd-11030;
parameter WEIGHT_0_3694 = 16'd4253;
parameter WEIGHT_0_3695 = 16'd2397;
parameter WEIGHT_0_3696 = 16'd3436;
parameter WEIGHT_0_3697 = 16'd4744;
parameter WEIGHT_0_3698 = 16'd-315;
parameter WEIGHT_0_3699 = 16'd8441;
parameter WEIGHT_0_3700 = 16'd2857;
parameter WEIGHT_0_3701 = 16'd-5708;
parameter WEIGHT_0_3702 = 16'd-21718;
parameter WEIGHT_0_3703 = 16'd-11366;
parameter WEIGHT_0_3704 = 16'd6543;
parameter WEIGHT_0_3705 = 16'd551;
parameter WEIGHT_0_3706 = 16'd8061;
parameter WEIGHT_0_3707 = 16'd1848;
parameter WEIGHT_0_3708 = 16'd-1060;
parameter WEIGHT_0_3709 = 16'd3495;
parameter WEIGHT_0_3710 = 16'd5547;
parameter WEIGHT_0_3711 = 16'd-4087;
parameter WEIGHT_0_3712 = 16'd-21101;
parameter WEIGHT_0_3713 = 16'd-13271;
parameter WEIGHT_0_3714 = 16'd6911;
parameter WEIGHT_0_3715 = 16'd2166;
parameter WEIGHT_0_3716 = 16'd4121;
parameter WEIGHT_0_3717 = 16'd567;
parameter WEIGHT_0_3718 = 16'd-4667;
parameter WEIGHT_0_3719 = 16'd3169;
parameter WEIGHT_0_3720 = 16'd1897;
parameter WEIGHT_0_3721 = 16'd-1316;
parameter WEIGHT_0_3722 = 16'd-14177;
parameter WEIGHT_0_3723 = 16'd-6372;
parameter WEIGHT_0_3724 = 16'd9195;
parameter WEIGHT_0_3725 = 16'd2050;
parameter WEIGHT_0_3726 = 16'd4293;
parameter WEIGHT_0_3727 = 16'd1351;
parameter WEIGHT_0_3728 = 16'd-4970;
parameter WEIGHT_0_3729 = 16'd3506;
parameter WEIGHT_0_3730 = 16'd3051;
parameter WEIGHT_0_3731 = 16'd-5149;
parameter WEIGHT_0_3732 = 16'd-8179;
parameter WEIGHT_0_3733 = 16'd-4554;
parameter WEIGHT_0_3734 = 16'd8086;
parameter WEIGHT_0_3735 = 16'd636;
parameter WEIGHT_0_3736 = 16'd3268;
parameter WEIGHT_0_3737 = 16'd-2853;
parameter WEIGHT_0_3738 = 16'd-2263;
parameter WEIGHT_0_3739 = 16'd3738;
parameter WEIGHT_0_3740 = 16'd324;
parameter WEIGHT_0_3741 = 16'd-16457;
parameter WEIGHT_0_3742 = 16'd-10166;
parameter WEIGHT_0_3743 = 16'd-4883;
parameter WEIGHT_0_3744 = 16'd11962;
parameter WEIGHT_0_3745 = 16'd6048;
parameter WEIGHT_0_3746 = 16'd3151;
parameter WEIGHT_0_3747 = 16'd-8061;
parameter WEIGHT_0_3748 = 16'd-8325;
parameter WEIGHT_0_3749 = 16'd-771;
parameter WEIGHT_0_3750 = 16'd150;
parameter WEIGHT_0_3751 = 16'd-14429;
parameter WEIGHT_0_3752 = 16'd-4688;
parameter WEIGHT_0_3753 = 16'd-3505;
parameter WEIGHT_0_3754 = 16'd15684;
parameter WEIGHT_0_3755 = 16'd8125;
parameter WEIGHT_0_3756 = 16'd2535;
parameter WEIGHT_0_3757 = 16'd-16183;
parameter WEIGHT_0_3758 = 16'd313;
parameter WEIGHT_0_3759 = 16'd-3694;
parameter WEIGHT_0_3760 = 16'd-744;
parameter WEIGHT_0_3761 = 16'd-8384;
parameter WEIGHT_0_3762 = 16'd-6042;
parameter WEIGHT_0_3763 = 16'd1956;
parameter WEIGHT_0_3764 = 16'd11193;
parameter WEIGHT_0_3765 = 16'd8730;
parameter WEIGHT_0_3766 = 16'd5341;
parameter WEIGHT_0_3767 = 16'd-24054;
parameter WEIGHT_0_3768 = 16'd4965;
parameter WEIGHT_0_3769 = 16'd-2951;
parameter WEIGHT_0_3770 = 16'd-13825;
parameter WEIGHT_0_3771 = 16'd10763;
parameter WEIGHT_0_3772 = 16'd-6544;
parameter WEIGHT_0_3773 = 16'd4479;
parameter WEIGHT_0_3774 = 16'd-2708;
parameter WEIGHT_0_3775 = 16'd5581;
parameter WEIGHT_0_3776 = 16'd-4853;
parameter WEIGHT_0_3777 = 16'd-26113;
parameter WEIGHT_0_3778 = 16'd7594;
parameter WEIGHT_0_3779 = 16'd-92;
parameter WEIGHT_0_3780 = 16'd-21460;
parameter WEIGHT_0_3781 = 16'd17480;
parameter WEIGHT_0_3782 = 16'd-6925;
parameter WEIGHT_0_3783 = 16'd3004;
parameter WEIGHT_0_3784 = 16'd-3214;
parameter WEIGHT_0_3785 = 16'd-2077;
parameter WEIGHT_0_3786 = 16'd-4934;
parameter WEIGHT_0_3787 = 16'd-11515;
parameter WEIGHT_0_3788 = 16'd3022;
parameter WEIGHT_0_3789 = 16'd6072;
parameter WEIGHT_0_3790 = 16'd-20627;
parameter WEIGHT_0_3791 = 16'd13751;
parameter WEIGHT_0_3792 = 16'd-6534;
parameter WEIGHT_0_3793 = 16'd1544;
parameter WEIGHT_0_3794 = 16'd1801;
parameter WEIGHT_0_3795 = 16'd-6401;
parameter WEIGHT_0_3796 = 16'd131;
parameter WEIGHT_0_3797 = 16'd312;
parameter WEIGHT_0_3798 = 16'd4654;
parameter WEIGHT_0_3799 = 16'd6308;
parameter WEIGHT_0_3800 = 16'd-18442;
parameter WEIGHT_0_3801 = 16'd2692;
parameter WEIGHT_0_3802 = 16'd-8084;
parameter WEIGHT_0_3803 = 16'd1182;
parameter WEIGHT_0_3804 = 16'd5903;
parameter WEIGHT_0_3805 = 16'd-13656;
parameter WEIGHT_0_3806 = 16'd-98;
parameter WEIGHT_0_3807 = 16'd2659;
parameter WEIGHT_0_3808 = 16'd461;
parameter WEIGHT_0_3809 = 16'd7749;
parameter WEIGHT_0_3810 = 16'd-8898;
parameter WEIGHT_0_3811 = 16'd-557;
parameter WEIGHT_0_3812 = 16'd-6480;
parameter WEIGHT_0_3813 = 16'd354;
parameter WEIGHT_0_3814 = 16'd7879;
parameter WEIGHT_0_3815 = 16'd-7243;
parameter WEIGHT_0_3816 = 16'd-2668;
parameter WEIGHT_0_3817 = 16'd5891;
parameter WEIGHT_0_3818 = 16'd-2495;
parameter WEIGHT_0_3819 = 16'd10204;
parameter WEIGHT_0_3820 = 16'd-248;
parameter WEIGHT_0_3821 = 16'd-5034;
parameter WEIGHT_0_3822 = 16'd-1810;
parameter WEIGHT_0_3823 = 16'd2344;
parameter WEIGHT_0_3824 = 16'd6437;
parameter WEIGHT_0_3825 = 16'd-7450;
parameter WEIGHT_0_3826 = 16'd-5841;
parameter WEIGHT_0_3827 = 16'd2005;
parameter WEIGHT_0_3828 = 16'd-2747;
parameter WEIGHT_0_3829 = 16'd7530;
parameter WEIGHT_0_3830 = 16'd-4572;
parameter WEIGHT_0_3831 = 16'd-10537;
parameter WEIGHT_0_3832 = 16'd-4568;
parameter WEIGHT_0_3833 = 16'd-2508;
parameter WEIGHT_0_3834 = 16'd5172;
parameter WEIGHT_0_3835 = 16'd-4829;
parameter WEIGHT_0_3836 = 16'd-1706;
parameter WEIGHT_0_3837 = 16'd1593;
parameter WEIGHT_0_3838 = 16'd1093;
parameter WEIGHT_0_3839 = 16'd9694;
parameter WEIGHT_0_3840 = 16'd-542;
parameter WEIGHT_0_3841 = 16'd-9712;
parameter WEIGHT_0_3842 = 16'd-4025;
parameter WEIGHT_0_3843 = 16'd-9689;
parameter WEIGHT_0_3844 = 16'd5362;
parameter WEIGHT_0_3845 = 16'd-5568;
parameter WEIGHT_0_3846 = 16'd-91;
parameter WEIGHT_0_3847 = 16'd1871;
parameter WEIGHT_0_3848 = 16'd2701;
parameter WEIGHT_0_3849 = 16'd6788;
parameter WEIGHT_0_3850 = 16'd1288;
parameter WEIGHT_0_3851 = 16'd-3918;
parameter WEIGHT_0_3852 = 16'd-2386;
parameter WEIGHT_0_3853 = 16'd-10623;
parameter WEIGHT_0_3854 = 16'd2871;
parameter WEIGHT_0_3855 = 16'd-10738;
parameter WEIGHT_0_3856 = 16'd2263;
parameter WEIGHT_0_3857 = 16'd-1351;
parameter WEIGHT_0_3858 = 16'd755;
parameter WEIGHT_0_3859 = 16'd5687;
parameter WEIGHT_0_3860 = 16'd4315;
parameter WEIGHT_0_3861 = 16'd-7954;
parameter WEIGHT_0_3862 = 16'd-8997;
parameter WEIGHT_0_3863 = 16'd-15684;
parameter WEIGHT_0_3864 = 16'd3289;
parameter WEIGHT_0_3865 = 16'd-11574;
parameter WEIGHT_0_3866 = 16'd8822;
parameter WEIGHT_0_3867 = 16'd1201;
parameter WEIGHT_0_3868 = 16'd-1257;
parameter WEIGHT_0_3869 = 16'd3581;
parameter WEIGHT_0_3870 = 16'd10639;
parameter WEIGHT_0_3871 = 16'd-14452;
parameter WEIGHT_0_3872 = 16'd-3960;
parameter WEIGHT_0_3873 = 16'd-11559;
parameter WEIGHT_0_3874 = 16'd-5144;
parameter WEIGHT_0_3875 = 16'd-21551;
parameter WEIGHT_0_3876 = 16'd10814;
parameter WEIGHT_0_3877 = 16'd-4581;
parameter WEIGHT_0_3878 = 16'd4315;
parameter WEIGHT_0_3879 = 16'd-7146;
parameter WEIGHT_0_3880 = 16'd6542;
parameter WEIGHT_0_3881 = 16'd-15180;
parameter WEIGHT_0_3882 = 16'd3050;
parameter WEIGHT_0_3883 = 16'd-7567;
parameter WEIGHT_0_3884 = 16'd-7256;
parameter WEIGHT_0_3885 = 16'd-18493;
parameter WEIGHT_0_3886 = 16'd7914;
parameter WEIGHT_0_3887 = 16'd-4875;
parameter WEIGHT_0_3888 = 16'd-484;
parameter WEIGHT_0_3889 = 16'd-16109;
parameter WEIGHT_0_3890 = 16'd-1019;
parameter WEIGHT_0_3891 = 16'd-6519;
parameter WEIGHT_0_3892 = 16'd12810;
parameter WEIGHT_0_3893 = 16'd-4519;
parameter WEIGHT_0_3894 = 16'd-1239;
parameter WEIGHT_0_3895 = 16'd-8706;
parameter WEIGHT_0_3896 = 16'd-4955;
parameter WEIGHT_0_3897 = 16'd-2632;
parameter WEIGHT_0_3898 = 16'd2888;
parameter WEIGHT_0_3899 = 16'd-16004;
parameter WEIGHT_0_3900 = 16'd-8725;
parameter WEIGHT_0_3901 = 16'd-5599;
parameter WEIGHT_0_3902 = 16'd15032;
parameter WEIGHT_0_3903 = 16'd-2969;
parameter WEIGHT_0_3904 = 16'd-4156;
parameter WEIGHT_0_3905 = 16'd-2158;
parameter WEIGHT_0_3906 = 16'd-13141;
parameter WEIGHT_0_3907 = 16'd-4440;
parameter WEIGHT_0_3908 = 16'd-3376;
parameter WEIGHT_0_3909 = 16'd-11068;
parameter WEIGHT_0_3910 = 16'd-2824;
parameter WEIGHT_0_3911 = 16'd-803;
parameter WEIGHT_0_3912 = 16'd4748;
parameter WEIGHT_0_3913 = 16'd-4200;
parameter WEIGHT_0_3914 = 16'd-4181;
parameter WEIGHT_0_3915 = 16'd-2008;
parameter WEIGHT_0_3916 = 16'd-7702;
parameter WEIGHT_0_3917 = 16'd-4616;
parameter WEIGHT_0_3918 = 16'd-1403;
parameter WEIGHT_0_3919 = 16'd-3242;
parameter WEIGHT_0_3920 = 16'd-1120;
parameter WEIGHT_0_3921 = 16'd782;
parameter WEIGHT_0_3922 = 16'd922;
parameter WEIGHT_0_3923 = 16'd-2772;
parameter WEIGHT_0_3924 = 16'd862;
parameter WEIGHT_0_3925 = 16'd4880;
parameter WEIGHT_0_3926 = 16'd-3024;
parameter WEIGHT_0_3927 = 16'd-3027;
parameter WEIGHT_0_3928 = 16'd-2107;
parameter WEIGHT_0_3929 = 16'd-2984;
parameter WEIGHT_0_3930 = 16'd-1631;
parameter WEIGHT_0_3931 = 16'd-2621;
parameter WEIGHT_0_3932 = 16'd-909;
parameter WEIGHT_0_3933 = 16'd5035;
parameter WEIGHT_0_3934 = 16'd-1046;
parameter WEIGHT_0_3935 = 16'd-2982;
parameter WEIGHT_0_3936 = 16'd-1304;
parameter WEIGHT_0_3937 = 16'd784;
parameter WEIGHT_0_3938 = 16'd-1494;
parameter WEIGHT_0_3939 = 16'd-1107;
parameter WEIGHT_0_3940 = 16'd-2503;
parameter WEIGHT_0_3941 = 16'd3257;
parameter WEIGHT_0_3942 = 16'd-932;
parameter WEIGHT_0_3943 = 16'd1756;
parameter WEIGHT_0_3944 = 16'd-5680;
parameter WEIGHT_0_3945 = 16'd-6142;
parameter WEIGHT_0_3946 = 16'd1196;
parameter WEIGHT_0_3947 = 16'd9102;
parameter WEIGHT_0_3948 = 16'd-7857;
parameter WEIGHT_0_3949 = 16'd-10813;
parameter WEIGHT_0_3950 = 16'd-10573;
parameter WEIGHT_0_3951 = 16'd4378;
parameter WEIGHT_0_3952 = 16'd-5212;
parameter WEIGHT_0_3953 = 16'd2679;
parameter WEIGHT_0_3954 = 16'd-2424;
parameter WEIGHT_0_3955 = 16'd-1668;
parameter WEIGHT_0_3956 = 16'd-10824;
parameter WEIGHT_0_3957 = 16'd7231;
parameter WEIGHT_0_3958 = 16'd-5944;
parameter WEIGHT_0_3959 = 16'd1780;
parameter WEIGHT_0_3960 = 16'd-6607;
parameter WEIGHT_0_3961 = 16'd4102;
parameter WEIGHT_0_3962 = 16'd-10325;
parameter WEIGHT_0_3963 = 16'd-3874;
parameter WEIGHT_0_3964 = 16'd4862;
parameter WEIGHT_0_3965 = 16'd-558;
parameter WEIGHT_0_3966 = 16'd-15097;
parameter WEIGHT_0_3967 = 16'd5399;
parameter WEIGHT_0_3968 = 16'd-13645;
parameter WEIGHT_0_3969 = 16'd4917;
parameter WEIGHT_0_3970 = 16'd5043;
parameter WEIGHT_0_3971 = 16'd-1719;
parameter WEIGHT_0_3972 = 16'd-12645;
parameter WEIGHT_0_3973 = 16'd-10365;
parameter WEIGHT_0_3974 = 16'd7845;
parameter WEIGHT_0_3975 = 16'd1094;
parameter WEIGHT_0_3976 = 16'd-300;
parameter WEIGHT_0_3977 = 16'd2004;
parameter WEIGHT_0_3978 = 16'd-5027;
parameter WEIGHT_0_3979 = 16'd3601;
parameter WEIGHT_0_3980 = 16'd6077;
parameter WEIGHT_0_3981 = 16'd-7466;
parameter WEIGHT_0_3982 = 16'd-12095;
parameter WEIGHT_0_3983 = 16'd-10545;
parameter WEIGHT_0_3984 = 16'd7388;
parameter WEIGHT_0_3985 = 16'd-3072;
parameter WEIGHT_0_3986 = 16'd1492;
parameter WEIGHT_0_3987 = 16'd-2619;
parameter WEIGHT_0_3988 = 16'd-8474;
parameter WEIGHT_0_3989 = 16'd2637;
parameter WEIGHT_0_3990 = 16'd4472;
parameter WEIGHT_0_3991 = 16'd-6364;
parameter WEIGHT_0_3992 = 16'd-6761;
parameter WEIGHT_0_3993 = 16'd-9546;
parameter WEIGHT_0_3994 = 16'd10279;
parameter WEIGHT_0_3995 = 16'd-952;
parameter WEIGHT_0_3996 = 16'd1043;
parameter WEIGHT_0_3997 = 16'd-3227;
parameter WEIGHT_0_3998 = 16'd-8939;
parameter WEIGHT_0_3999 = 16'd3452;
parameter WEIGHT_0_4000 = 16'd2517;
parameter WEIGHT_0_4001 = 16'd-502;
parameter WEIGHT_0_4002 = 16'd-2787;
parameter WEIGHT_0_4003 = 16'd-4142;
parameter WEIGHT_0_4004 = 16'd8976;
parameter WEIGHT_0_4005 = 16'd-699;
parameter WEIGHT_0_4006 = 16'd2331;
parameter WEIGHT_0_4007 = 16'd-3916;
parameter WEIGHT_0_4008 = 16'd-5325;
parameter WEIGHT_0_4009 = 16'd4019;
parameter WEIGHT_0_4010 = 16'd1880;
parameter WEIGHT_0_4011 = 16'd-6970;
parameter WEIGHT_0_4012 = 16'd-3370;
parameter WEIGHT_0_4013 = 16'd-6300;
parameter WEIGHT_0_4014 = 16'd8576;
parameter WEIGHT_0_4015 = 16'd4538;
parameter WEIGHT_0_4016 = 16'd3271;
parameter WEIGHT_0_4017 = 16'd-6780;
parameter WEIGHT_0_4018 = 16'd-9056;
parameter WEIGHT_0_4019 = 16'd-694;
parameter WEIGHT_0_4020 = 16'd3798;
parameter WEIGHT_0_4021 = 16'd-17449;
parameter WEIGHT_0_4022 = 16'd-1328;
parameter WEIGHT_0_4023 = 16'd-6575;
parameter WEIGHT_0_4024 = 16'd7918;
parameter WEIGHT_0_4025 = 16'd3967;
parameter WEIGHT_0_4026 = 16'd6556;
parameter WEIGHT_0_4027 = 16'd-9277;
parameter WEIGHT_0_4028 = 16'd-2590;
parameter WEIGHT_0_4029 = 16'd20;
parameter WEIGHT_0_4030 = 16'd4231;
parameter WEIGHT_0_4031 = 16'd-17664;
parameter WEIGHT_0_4032 = 16'd-1702;
parameter WEIGHT_0_4033 = 16'd-4758;
parameter WEIGHT_0_4034 = 16'd9800;
parameter WEIGHT_0_4035 = 16'd4502;
parameter WEIGHT_0_4036 = 16'd5445;
parameter WEIGHT_0_4037 = 16'd-19242;
parameter WEIGHT_0_4038 = 16'd951;
parameter WEIGHT_0_4039 = 16'd-3718;
parameter WEIGHT_0_4040 = 16'd-4282;
parameter WEIGHT_0_4041 = 16'd-5085;
parameter WEIGHT_0_4042 = 16'd1090;
parameter WEIGHT_0_4043 = 16'd2275;
parameter WEIGHT_0_4044 = 16'd3839;
parameter WEIGHT_0_4045 = 16'd2294;
parameter WEIGHT_0_4046 = 16'd4366;
parameter WEIGHT_0_4047 = 16'd-26662;
parameter WEIGHT_0_4048 = 16'd6123;
parameter WEIGHT_0_4049 = 16'd-3903;
parameter WEIGHT_0_4050 = 16'd-10145;
parameter WEIGHT_0_4051 = 16'd9552;
parameter WEIGHT_0_4052 = 16'd4631;
parameter WEIGHT_0_4053 = 16'd2202;
parameter WEIGHT_0_4054 = 16'd-3445;
parameter WEIGHT_0_4055 = 16'd1346;
parameter WEIGHT_0_4056 = 16'd124;
parameter WEIGHT_0_4057 = 16'd-16786;
parameter WEIGHT_0_4058 = 16'd9162;
parameter WEIGHT_0_4059 = 16'd1497;
parameter WEIGHT_0_4060 = 16'd-23183;
parameter WEIGHT_0_4061 = 16'd13273;
parameter WEIGHT_0_4062 = 16'd-458;
parameter WEIGHT_0_4063 = 16'd3215;
parameter WEIGHT_0_4064 = 16'd-124;
parameter WEIGHT_0_4065 = 16'd-3958;
parameter WEIGHT_0_4066 = 16'd-1004;
parameter WEIGHT_0_4067 = 16'd-7488;
parameter WEIGHT_0_4068 = 16'd4705;
parameter WEIGHT_0_4069 = 16'd-384;
parameter WEIGHT_0_4070 = 16'd-19164;
parameter WEIGHT_0_4071 = 16'd11278;
parameter WEIGHT_0_4072 = 16'd-2147;
parameter WEIGHT_0_4073 = 16'd-1400;
parameter WEIGHT_0_4074 = 16'd4467;
parameter WEIGHT_0_4075 = 16'd-5053;
parameter WEIGHT_0_4076 = 16'd164;
parameter WEIGHT_0_4077 = 16'd-3483;
parameter WEIGHT_0_4078 = 16'd1331;
parameter WEIGHT_0_4079 = 16'd5210;
parameter WEIGHT_0_4080 = 16'd-19097;
parameter WEIGHT_0_4081 = 16'd-1391;
parameter WEIGHT_0_4082 = 16'd-4509;
parameter WEIGHT_0_4083 = 16'd272;
parameter WEIGHT_0_4084 = 16'd8728;
parameter WEIGHT_0_4085 = 16'd-10160;
parameter WEIGHT_0_4086 = 16'd2292;
parameter WEIGHT_0_4087 = 16'd443;
parameter WEIGHT_0_4088 = 16'd430;
parameter WEIGHT_0_4089 = 16'd7547;
parameter WEIGHT_0_4090 = 16'd-8541;
parameter WEIGHT_0_4091 = 16'd-8710;
parameter WEIGHT_0_4092 = 16'd-6708;
parameter WEIGHT_0_4093 = 16'd-748;
parameter WEIGHT_0_4094 = 16'd11276;
parameter WEIGHT_0_4095 = 16'd-6000;
parameter WEIGHT_0_4096 = 16'd-6182;
parameter WEIGHT_0_4097 = 16'd4473;
parameter WEIGHT_0_4098 = 16'd-1578;
parameter WEIGHT_0_4099 = 16'd8249;
parameter WEIGHT_0_4100 = 16'd-3154;
parameter WEIGHT_0_4101 = 16'd-11489;
parameter WEIGHT_0_4102 = 16'd-4501;
parameter WEIGHT_0_4103 = 16'd1277;
parameter WEIGHT_0_4104 = 16'd8095;
parameter WEIGHT_0_4105 = 16'd-6246;
parameter WEIGHT_0_4106 = 16'd-4796;
parameter WEIGHT_0_4107 = 16'd8202;
parameter WEIGHT_0_4108 = 16'd-4844;
parameter WEIGHT_0_4109 = 16'd4294;
parameter WEIGHT_0_4110 = 16'd-4034;
parameter WEIGHT_0_4111 = 16'd-12119;
parameter WEIGHT_0_4112 = 16'd-4806;
parameter WEIGHT_0_4113 = 16'd-2183;
parameter WEIGHT_0_4114 = 16'd5350;
parameter WEIGHT_0_4115 = 16'd-3033;
parameter WEIGHT_0_4116 = 16'd-2257;
parameter WEIGHT_0_4117 = 16'd6439;
parameter WEIGHT_0_4118 = 16'd-4120;
parameter WEIGHT_0_4119 = 16'd3862;
parameter WEIGHT_0_4120 = 16'd197;
parameter WEIGHT_0_4121 = 16'd-7552;
parameter WEIGHT_0_4122 = 16'd-2527;
parameter WEIGHT_0_4123 = 16'd-5083;
parameter WEIGHT_0_4124 = 16'd6344;
parameter WEIGHT_0_4125 = 16'd146;
parameter WEIGHT_0_4126 = 16'd2529;
parameter WEIGHT_0_4127 = 16'd8089;
parameter WEIGHT_0_4128 = 16'd-5466;
parameter WEIGHT_0_4129 = 16'd1776;
parameter WEIGHT_0_4130 = 16'd3917;
parameter WEIGHT_0_4131 = 16'd-8255;
parameter WEIGHT_0_4132 = 16'd-3649;
parameter WEIGHT_0_4133 = 16'd-1639;
parameter WEIGHT_0_4134 = 16'd3129;
parameter WEIGHT_0_4135 = 16'd-3300;
parameter WEIGHT_0_4136 = 16'd3105;
parameter WEIGHT_0_4137 = 16'd2392;
parameter WEIGHT_0_4138 = 16'd-8346;
parameter WEIGHT_0_4139 = 16'd2499;
parameter WEIGHT_0_4140 = 16'd5152;
parameter WEIGHT_0_4141 = 16'd-8019;
parameter WEIGHT_0_4142 = 16'd-6647;
parameter WEIGHT_0_4143 = 16'd-6313;
parameter WEIGHT_0_4144 = 16'd-681;
parameter WEIGHT_0_4145 = 16'd-2883;
parameter WEIGHT_0_4146 = 16'd5669;
parameter WEIGHT_0_4147 = 16'd4161;
parameter WEIGHT_0_4148 = 16'd-9212;
parameter WEIGHT_0_4149 = 16'd-4912;
parameter WEIGHT_0_4150 = 16'd7000;
parameter WEIGHT_0_4151 = 16'd-8356;
parameter WEIGHT_0_4152 = 16'd-3405;
parameter WEIGHT_0_4153 = 16'd-5593;
parameter WEIGHT_0_4154 = 16'd-4050;
parameter WEIGHT_0_4155 = 16'd-5257;
parameter WEIGHT_0_4156 = 16'd10426;
parameter WEIGHT_0_4157 = 16'd4119;
parameter WEIGHT_0_4158 = 16'd-8709;
parameter WEIGHT_0_4159 = 16'd-9608;
parameter WEIGHT_0_4160 = 16'd10087;
parameter WEIGHT_0_4161 = 16'd-7431;
parameter WEIGHT_0_4162 = 16'd2730;
parameter WEIGHT_0_4163 = 16'd-6985;
parameter WEIGHT_0_4164 = 16'd-5311;
parameter WEIGHT_0_4165 = 16'd-6428;
parameter WEIGHT_0_4166 = 16'd6132;
parameter WEIGHT_0_4167 = 16'd-1440;
parameter WEIGHT_0_4168 = 16'd-8897;
parameter WEIGHT_0_4169 = 16'd-20760;
parameter WEIGHT_0_4170 = 16'd1853;
parameter WEIGHT_0_4171 = 16'd-5646;
parameter WEIGHT_0_4172 = 16'd12392;
parameter WEIGHT_0_4173 = 16'd-11044;
parameter WEIGHT_0_4174 = 16'd-7854;
parameter WEIGHT_0_4175 = 16'd-11740;
parameter WEIGHT_0_4176 = 16'd-2300;
parameter WEIGHT_0_4177 = 16'd-3710;
parameter WEIGHT_0_4178 = 16'd-1146;
parameter WEIGHT_0_4179 = 16'd-14937;
parameter WEIGHT_0_4180 = 16'd-11345;
parameter WEIGHT_0_4181 = 16'd-3670;
parameter WEIGHT_0_4182 = 16'd13069;
parameter WEIGHT_0_4183 = 16'd-7486;
parameter WEIGHT_0_4184 = 16'd-7308;
parameter WEIGHT_0_4185 = 16'd-9016;
parameter WEIGHT_0_4186 = 16'd-9719;
parameter WEIGHT_0_4187 = 16'd-6059;
parameter WEIGHT_0_4188 = 16'd-10671;
parameter WEIGHT_0_4189 = 16'd-8871;
parameter WEIGHT_0_4190 = 16'd-4856;
parameter WEIGHT_0_4191 = 16'd-1505;
parameter WEIGHT_0_4192 = 16'd6771;
parameter WEIGHT_0_4193 = 16'd-5169;
parameter WEIGHT_0_4194 = 16'd-4749;
parameter WEIGHT_0_4195 = 16'd-4125;
parameter WEIGHT_0_4196 = 16'd-3038;
parameter WEIGHT_0_4197 = 16'd-5628;
parameter WEIGHT_0_4198 = 16'd-6698;
parameter WEIGHT_0_4199 = 16'd-6858;
parameter WEIGHT_0_4200 = 16'd-3713;
parameter WEIGHT_0_4201 = 16'd1629;
parameter WEIGHT_0_4202 = 16'd18;
parameter WEIGHT_0_4203 = 16'd-273;
parameter WEIGHT_0_4204 = 16'd-3998;
parameter WEIGHT_0_4205 = 16'd878;
parameter WEIGHT_0_4206 = 16'd-2952;
parameter WEIGHT_0_4207 = 16'd-1204;
parameter WEIGHT_0_4208 = 16'd-3211;
parameter WEIGHT_0_4209 = 16'd277;
parameter WEIGHT_0_4210 = 16'd-3722;
parameter WEIGHT_0_4211 = 16'd-254;
parameter WEIGHT_0_4212 = 16'd-3656;
parameter WEIGHT_0_4213 = 16'd4506;
parameter WEIGHT_0_4214 = 16'd1905;
parameter WEIGHT_0_4215 = 16'd-5033;
parameter WEIGHT_0_4216 = 16'd-2608;
parameter WEIGHT_0_4217 = 16'd-3653;
parameter WEIGHT_0_4218 = 16'd-3895;
parameter WEIGHT_0_4219 = 16'd861;
parameter WEIGHT_0_4220 = 16'd-3562;
parameter WEIGHT_0_4221 = 16'd585;
parameter WEIGHT_0_4222 = 16'd-2750;
parameter WEIGHT_0_4223 = 16'd3502;
parameter WEIGHT_0_4224 = 16'd3401;
parameter WEIGHT_0_4225 = 16'd-7705;
parameter WEIGHT_0_4226 = 16'd-4830;
parameter WEIGHT_0_4227 = 16'd2648;
parameter WEIGHT_0_4228 = 16'd-10254;
parameter WEIGHT_0_4229 = 16'd-7080;
parameter WEIGHT_0_4230 = 16'd-11432;
parameter WEIGHT_0_4231 = 16'd1183;
parameter WEIGHT_0_4232 = 16'd741;
parameter WEIGHT_0_4233 = 16'd2218;
parameter WEIGHT_0_4234 = 16'd1189;
parameter WEIGHT_0_4235 = 16'd-2218;
parameter WEIGHT_0_4236 = 16'd-13132;
parameter WEIGHT_0_4237 = 16'd4123;
parameter WEIGHT_0_4238 = 16'd-6974;
parameter WEIGHT_0_4239 = 16'd-1234;
parameter WEIGHT_0_4240 = 16'd1194;
parameter WEIGHT_0_4241 = 16'd-3697;
parameter WEIGHT_0_4242 = 16'd-1383;
parameter WEIGHT_0_4243 = 16'd-2091;
parameter WEIGHT_0_4244 = 16'd5497;
parameter WEIGHT_0_4245 = 16'd-6221;
parameter WEIGHT_0_4246 = 16'd-19270;
parameter WEIGHT_0_4247 = 16'd1024;
parameter WEIGHT_0_4248 = 16'd-13487;
parameter WEIGHT_0_4249 = 16'd1974;
parameter WEIGHT_0_4250 = 16'd3672;
parameter WEIGHT_0_4251 = 16'd-9704;
parameter WEIGHT_0_4252 = 16'd1734;
parameter WEIGHT_0_4253 = 16'd-1938;
parameter WEIGHT_0_4254 = 16'd2248;
parameter WEIGHT_0_4255 = 16'd-8170;
parameter WEIGHT_0_4256 = 16'd-204;
parameter WEIGHT_0_4257 = 16'd814;
parameter WEIGHT_0_4258 = 16'd-11177;
parameter WEIGHT_0_4259 = 16'd2213;
parameter WEIGHT_0_4260 = 16'd1735;
parameter WEIGHT_0_4261 = 16'd-9831;
parameter WEIGHT_0_4262 = 16'd-866;
parameter WEIGHT_0_4263 = 16'd-6033;
parameter WEIGHT_0_4264 = 16'd6039;
parameter WEIGHT_0_4265 = 16'd-4655;
parameter WEIGHT_0_4266 = 16'd2842;
parameter WEIGHT_0_4267 = 16'd18;
parameter WEIGHT_0_4268 = 16'd-9318;
parameter WEIGHT_0_4269 = 16'd-1383;
parameter WEIGHT_0_4270 = 16'd8076;
parameter WEIGHT_0_4271 = 16'd-7586;
parameter WEIGHT_0_4272 = 16'd-852;
parameter WEIGHT_0_4273 = 16'd-11771;
parameter WEIGHT_0_4274 = 16'd6103;
parameter WEIGHT_0_4275 = 16'd-5873;
parameter WEIGHT_0_4276 = 16'd5383;
parameter WEIGHT_0_4277 = 16'd-3203;
parameter WEIGHT_0_4278 = 16'd-8058;
parameter WEIGHT_0_4279 = 16'd2099;
parameter WEIGHT_0_4280 = 16'd6316;
parameter WEIGHT_0_4281 = 16'd-3403;
parameter WEIGHT_0_4282 = 16'd-1425;
parameter WEIGHT_0_4283 = 16'd-9868;
parameter WEIGHT_0_4284 = 16'd8690;
parameter WEIGHT_0_4285 = 16'd-2619;
parameter WEIGHT_0_4286 = 16'd4383;
parameter WEIGHT_0_4287 = 16'd-8231;
parameter WEIGHT_0_4288 = 16'd-7156;
parameter WEIGHT_0_4289 = 16'd-559;
parameter WEIGHT_0_4290 = 16'd3489;
parameter WEIGHT_0_4291 = 16'd-6873;
parameter WEIGHT_0_4292 = 16'd-2262;
parameter WEIGHT_0_4293 = 16'd-6562;
parameter WEIGHT_0_4294 = 16'd4391;
parameter WEIGHT_0_4295 = 16'd1837;
parameter WEIGHT_0_4296 = 16'd3870;
parameter WEIGHT_0_4297 = 16'd-8145;
parameter WEIGHT_0_4298 = 16'd-5308;
parameter WEIGHT_0_4299 = 16'd-2242;
parameter WEIGHT_0_4300 = 16'd5941;
parameter WEIGHT_0_4301 = 16'd-11340;
parameter WEIGHT_0_4302 = 16'd-56;
parameter WEIGHT_0_4303 = 16'd-5514;
parameter WEIGHT_0_4304 = 16'd7077;
parameter WEIGHT_0_4305 = 16'd2013;
parameter WEIGHT_0_4306 = 16'd9998;
parameter WEIGHT_0_4307 = 16'd-10549;
parameter WEIGHT_0_4308 = 16'd-3402;
parameter WEIGHT_0_4309 = 16'd721;
parameter WEIGHT_0_4310 = 16'd311;
parameter WEIGHT_0_4311 = 16'd-9046;
parameter WEIGHT_0_4312 = 16'd483;
parameter WEIGHT_0_4313 = 16'd-2844;
parameter WEIGHT_0_4314 = 16'd6593;
parameter WEIGHT_0_4315 = 16'd3636;
parameter WEIGHT_0_4316 = 16'd9217;
parameter WEIGHT_0_4317 = 16'd-15256;
parameter WEIGHT_0_4318 = 16'd1727;
parameter WEIGHT_0_4319 = 16'd-1572;
parameter WEIGHT_0_4320 = 16'd-4229;
parameter WEIGHT_0_4321 = 16'd535;
parameter WEIGHT_0_4322 = 16'd1239;
parameter WEIGHT_0_4323 = 16'd2546;
parameter WEIGHT_0_4324 = 16'd2943;
parameter WEIGHT_0_4325 = 16'd234;
parameter WEIGHT_0_4326 = 16'd1960;
parameter WEIGHT_0_4327 = 16'd-16946;
parameter WEIGHT_0_4328 = 16'd4457;
parameter WEIGHT_0_4329 = 16'd-2118;
parameter WEIGHT_0_4330 = 16'd-17717;
parameter WEIGHT_0_4331 = 16'd12256;
parameter WEIGHT_0_4332 = 16'd6477;
parameter WEIGHT_0_4333 = 16'd248;
parameter WEIGHT_0_4334 = 16'd-2595;
parameter WEIGHT_0_4335 = 16'd-608;
parameter WEIGHT_0_4336 = 16'd-205;
parameter WEIGHT_0_4337 = 16'd-12298;
parameter WEIGHT_0_4338 = 16'd8945;
parameter WEIGHT_0_4339 = 16'd-5134;
parameter WEIGHT_0_4340 = 16'd-23227;
parameter WEIGHT_0_4341 = 16'd16369;
parameter WEIGHT_0_4342 = 16'd-1608;
parameter WEIGHT_0_4343 = 16'd2811;
parameter WEIGHT_0_4344 = 16'd1675;
parameter WEIGHT_0_4345 = 16'd-9221;
parameter WEIGHT_0_4346 = 16'd1437;
parameter WEIGHT_0_4347 = 16'd-7687;
parameter WEIGHT_0_4348 = 16'd3642;
parameter WEIGHT_0_4349 = 16'd-2828;
parameter WEIGHT_0_4350 = 16'd-18640;
parameter WEIGHT_0_4351 = 16'd9232;
parameter WEIGHT_0_4352 = 16'd1340;
parameter WEIGHT_0_4353 = 16'd148;
parameter WEIGHT_0_4354 = 16'd8320;
parameter WEIGHT_0_4355 = 16'd-10173;
parameter WEIGHT_0_4356 = 16'd2346;
parameter WEIGHT_0_4357 = 16'd1122;
parameter WEIGHT_0_4358 = 16'd2032;
parameter WEIGHT_0_4359 = 16'd1096;
parameter WEIGHT_0_4360 = 16'd-16132;
parameter WEIGHT_0_4361 = 16'd-1113;
parameter WEIGHT_0_4362 = 16'd-2719;
parameter WEIGHT_0_4363 = 16'd-4309;
parameter WEIGHT_0_4364 = 16'd10249;
parameter WEIGHT_0_4365 = 16'd-8809;
parameter WEIGHT_0_4366 = 16'd-1095;
parameter WEIGHT_0_4367 = 16'd983;
parameter WEIGHT_0_4368 = 16'd-2032;
parameter WEIGHT_0_4369 = 16'd9370;
parameter WEIGHT_0_4370 = 16'd-4708;
parameter WEIGHT_0_4371 = 16'd-11226;
parameter WEIGHT_0_4372 = 16'd-548;
parameter WEIGHT_0_4373 = 16'd-621;
parameter WEIGHT_0_4374 = 16'd11473;
parameter WEIGHT_0_4375 = 16'd-4043;
parameter WEIGHT_0_4376 = 16'd-956;
parameter WEIGHT_0_4377 = 16'd7040;
parameter WEIGHT_0_4378 = 16'd-3595;
parameter WEIGHT_0_4379 = 16'd6891;
parameter WEIGHT_0_4380 = 16'd-2238;
parameter WEIGHT_0_4381 = 16'd-15520;
parameter WEIGHT_0_4382 = 16'd-3701;
parameter WEIGHT_0_4383 = 16'd-2356;
parameter WEIGHT_0_4384 = 16'd4303;
parameter WEIGHT_0_4385 = 16'd-2031;
parameter WEIGHT_0_4386 = 16'd-4344;
parameter WEIGHT_0_4387 = 16'd9532;
parameter WEIGHT_0_4388 = 16'd-3222;
parameter WEIGHT_0_4389 = 16'd-528;
parameter WEIGHT_0_4390 = 16'd-3527;
parameter WEIGHT_0_4391 = 16'd-16057;
parameter WEIGHT_0_4392 = 16'd-3692;
parameter WEIGHT_0_4393 = 16'd-4;
parameter WEIGHT_0_4394 = 16'd4480;
parameter WEIGHT_0_4395 = 16'd-3718;
parameter WEIGHT_0_4396 = 16'd411;
parameter WEIGHT_0_4397 = 16'd9817;
parameter WEIGHT_0_4398 = 16'd-7186;
parameter WEIGHT_0_4399 = 16'd-2028;
parameter WEIGHT_0_4400 = 16'd271;
parameter WEIGHT_0_4401 = 16'd-12408;
parameter WEIGHT_0_4402 = 16'd-5688;
parameter WEIGHT_0_4403 = 16'd3770;
parameter WEIGHT_0_4404 = 16'd233;
parameter WEIGHT_0_4405 = 16'd-5477;
parameter WEIGHT_0_4406 = 16'd390;
parameter WEIGHT_0_4407 = 16'd7822;
parameter WEIGHT_0_4408 = 16'd-9434;
parameter WEIGHT_0_4409 = 16'd-944;
parameter WEIGHT_0_4410 = 16'd2792;
parameter WEIGHT_0_4411 = 16'd-8404;
parameter WEIGHT_0_4412 = 16'd-7110;
parameter WEIGHT_0_4413 = 16'd3745;
parameter WEIGHT_0_4414 = 16'd-4062;
parameter WEIGHT_0_4415 = 16'd-932;
parameter WEIGHT_0_4416 = 16'd2089;
parameter WEIGHT_0_4417 = 16'd9469;
parameter WEIGHT_0_4418 = 16'd-7048;
parameter WEIGHT_0_4419 = 16'd-4951;
parameter WEIGHT_0_4420 = 16'd3726;
parameter WEIGHT_0_4421 = 16'd-10186;
parameter WEIGHT_0_4422 = 16'd-3938;
parameter WEIGHT_0_4423 = 16'd620;
parameter WEIGHT_0_4424 = 16'd166;
parameter WEIGHT_0_4425 = 16'd-1893;
parameter WEIGHT_0_4426 = 16'd4130;
parameter WEIGHT_0_4427 = 16'd6175;
parameter WEIGHT_0_4428 = 16'd-5839;
parameter WEIGHT_0_4429 = 16'd-3725;
parameter WEIGHT_0_4430 = 16'd4415;
parameter WEIGHT_0_4431 = 16'd-9705;
parameter WEIGHT_0_4432 = 16'd-1335;
parameter WEIGHT_0_4433 = 16'd3326;
parameter WEIGHT_0_4434 = 16'd-1534;
parameter WEIGHT_0_4435 = 16'd1411;
parameter WEIGHT_0_4436 = 16'd1617;
parameter WEIGHT_0_4437 = 16'd1415;
parameter WEIGHT_0_4438 = 16'd-9147;
parameter WEIGHT_0_4439 = 16'd-13307;
parameter WEIGHT_0_4440 = 16'd5167;
parameter WEIGHT_0_4441 = 16'd-12174;
parameter WEIGHT_0_4442 = 16'd7662;
parameter WEIGHT_0_4443 = 16'd2140;
parameter WEIGHT_0_4444 = 16'd-12908;
parameter WEIGHT_0_4445 = 16'd-692;
parameter WEIGHT_0_4446 = 16'd2313;
parameter WEIGHT_0_4447 = 16'd-1332;
parameter WEIGHT_0_4448 = 16'd-10151;
parameter WEIGHT_0_4449 = 16'd-21598;
parameter WEIGHT_0_4450 = 16'd-3349;
parameter WEIGHT_0_4451 = 16'd-5189;
parameter WEIGHT_0_4452 = 16'd13007;
parameter WEIGHT_0_4453 = 16'd-13250;
parameter WEIGHT_0_4454 = 16'd-7716;
parameter WEIGHT_0_4455 = 16'd-8725;
parameter WEIGHT_0_4456 = 16'd-2719;
parameter WEIGHT_0_4457 = 16'd-8363;
parameter WEIGHT_0_4458 = 16'd-5213;
parameter WEIGHT_0_4459 = 16'd-16831;
parameter WEIGHT_0_4460 = 16'd-11397;
parameter WEIGHT_0_4461 = 16'd-7807;
parameter WEIGHT_0_4462 = 16'd16028;
parameter WEIGHT_0_4463 = 16'd429;
parameter WEIGHT_0_4464 = 16'd-3958;
parameter WEIGHT_0_4465 = 16'd-12364;
parameter WEIGHT_0_4466 = 16'd-11196;
parameter WEIGHT_0_4467 = 16'd-5178;
parameter WEIGHT_0_4468 = 16'd-11097;
parameter WEIGHT_0_4469 = 16'd-5920;
parameter WEIGHT_0_4470 = 16'd-3814;
parameter WEIGHT_0_4471 = 16'd-6743;
parameter WEIGHT_0_4472 = 16'd5947;
parameter WEIGHT_0_4473 = 16'd-4994;
parameter WEIGHT_0_4474 = 16'd-877;
parameter WEIGHT_0_4475 = 16'd-4819;
parameter WEIGHT_0_4476 = 16'd-7875;
parameter WEIGHT_0_4477 = 16'd-3726;
parameter WEIGHT_0_4478 = 16'd-7724;
parameter WEIGHT_0_4479 = 16'd-3796;
parameter WEIGHT_0_4480 = 16'd194;
parameter WEIGHT_0_4481 = 16'd579;
parameter WEIGHT_0_4482 = 16'd-1943;
parameter WEIGHT_0_4483 = 16'd-3943;
parameter WEIGHT_0_4484 = 16'd-1984;
parameter WEIGHT_0_4485 = 16'd-186;
parameter WEIGHT_0_4486 = 16'd-2130;
parameter WEIGHT_0_4487 = 16'd4536;
parameter WEIGHT_0_4488 = 16'd248;
parameter WEIGHT_0_4489 = 16'd-3944;
parameter WEIGHT_0_4490 = 16'd-695;
parameter WEIGHT_0_4491 = 16'd5062;
parameter WEIGHT_0_4492 = 16'd-2800;
parameter WEIGHT_0_4493 = 16'd4884;
parameter WEIGHT_0_4494 = 16'd183;
parameter WEIGHT_0_4495 = 16'd-2995;
parameter WEIGHT_0_4496 = 16'd-11;
parameter WEIGHT_0_4497 = 16'd-2996;
parameter WEIGHT_0_4498 = 16'd-2738;
parameter WEIGHT_0_4499 = 16'd-4764;
parameter WEIGHT_0_4500 = 16'd-2099;
parameter WEIGHT_0_4501 = 16'd971;
parameter WEIGHT_0_4502 = 16'd-1182;
parameter WEIGHT_0_4503 = 16'd4336;
parameter WEIGHT_0_4504 = 16'd-488;
parameter WEIGHT_0_4505 = 16'd-9720;
parameter WEIGHT_0_4506 = 16'd-3855;
parameter WEIGHT_0_4507 = 16'd-2539;
parameter WEIGHT_0_4508 = 16'd-5887;
parameter WEIGHT_0_4509 = 16'd-9322;
parameter WEIGHT_0_4510 = 16'd-11190;
parameter WEIGHT_0_4511 = 16'd-1071;
parameter WEIGHT_0_4512 = 16'd4778;
parameter WEIGHT_0_4513 = 16'd4724;
parameter WEIGHT_0_4514 = 16'd-6387;
parameter WEIGHT_0_4515 = 16'd-89;
parameter WEIGHT_0_4516 = 16'd-10825;
parameter WEIGHT_0_4517 = 16'd-2323;
parameter WEIGHT_0_4518 = 16'd-6033;
parameter WEIGHT_0_4519 = 16'd-1769;
parameter WEIGHT_0_4520 = 16'd1285;
parameter WEIGHT_0_4521 = 16'd-7302;
parameter WEIGHT_0_4522 = 16'd4872;
parameter WEIGHT_0_4523 = 16'd3580;
parameter WEIGHT_0_4524 = 16'd-6586;
parameter WEIGHT_0_4525 = 16'd-1443;
parameter WEIGHT_0_4526 = 16'd-18997;
parameter WEIGHT_0_4527 = 16'd2774;
parameter WEIGHT_0_4528 = 16'd-14091;
parameter WEIGHT_0_4529 = 16'd2295;
parameter WEIGHT_0_4530 = 16'd7534;
parameter WEIGHT_0_4531 = 16'd-9419;
parameter WEIGHT_0_4532 = 16'd4699;
parameter WEIGHT_0_4533 = 16'd-183;
parameter WEIGHT_0_4534 = 16'd-2016;
parameter WEIGHT_0_4535 = 16'd-5754;
parameter WEIGHT_0_4536 = 16'd-1058;
parameter WEIGHT_0_4537 = 16'd-2099;
parameter WEIGHT_0_4538 = 16'd-14064;
parameter WEIGHT_0_4539 = 16'd882;
parameter WEIGHT_0_4540 = 16'd3782;
parameter WEIGHT_0_4541 = 16'd-12503;
parameter WEIGHT_0_4542 = 16'd5028;
parameter WEIGHT_0_4543 = 16'd-4626;
parameter WEIGHT_0_4544 = 16'd1428;
parameter WEIGHT_0_4545 = 16'd-5256;
parameter WEIGHT_0_4546 = 16'd810;
parameter WEIGHT_0_4547 = 16'd-1792;
parameter WEIGHT_0_4548 = 16'd-8761;
parameter WEIGHT_0_4549 = 16'd-703;
parameter WEIGHT_0_4550 = 16'd4063;
parameter WEIGHT_0_4551 = 16'd-9823;
parameter WEIGHT_0_4552 = 16'd-1111;
parameter WEIGHT_0_4553 = 16'd-5011;
parameter WEIGHT_0_4554 = 16'd5582;
parameter WEIGHT_0_4555 = 16'd-13492;
parameter WEIGHT_0_4556 = 16'd969;
parameter WEIGHT_0_4557 = 16'd2458;
parameter WEIGHT_0_4558 = 16'd-5102;
parameter WEIGHT_0_4559 = 16'd-418;
parameter WEIGHT_0_4560 = 16'd5053;
parameter WEIGHT_0_4561 = 16'd-9669;
parameter WEIGHT_0_4562 = 16'd-4177;
parameter WEIGHT_0_4563 = 16'd-11167;
parameter WEIGHT_0_4564 = 16'd10319;
parameter WEIGHT_0_4565 = 16'd-12561;
parameter WEIGHT_0_4566 = 16'd3741;
parameter WEIGHT_0_4567 = 16'd-4730;
parameter WEIGHT_0_4568 = 16'd-1257;
parameter WEIGHT_0_4569 = 16'd3868;
parameter WEIGHT_0_4570 = 16'd7349;
parameter WEIGHT_0_4571 = 16'd-7211;
parameter WEIGHT_0_4572 = 16'd349;
parameter WEIGHT_0_4573 = 16'd-11228;
parameter WEIGHT_0_4574 = 16'd5097;
parameter WEIGHT_0_4575 = 16'd-7280;
parameter WEIGHT_0_4576 = 16'd8276;
parameter WEIGHT_0_4577 = 16'd-9049;
parameter WEIGHT_0_4578 = 16'd1333;
parameter WEIGHT_0_4579 = 16'd-1279;
parameter WEIGHT_0_4580 = 16'd4213;
parameter WEIGHT_0_4581 = 16'd-2848;
parameter WEIGHT_0_4582 = 16'd3442;
parameter WEIGHT_0_4583 = 16'd-5922;
parameter WEIGHT_0_4584 = 16'd-1459;
parameter WEIGHT_0_4585 = 16'd-4772;
parameter WEIGHT_0_4586 = 16'd8961;
parameter WEIGHT_0_4587 = 16'd-9496;
parameter WEIGHT_0_4588 = 16'd-336;
parameter WEIGHT_0_4589 = 16'd985;
parameter WEIGHT_0_4590 = 16'd1907;
parameter WEIGHT_0_4591 = 16'd-6874;
parameter WEIGHT_0_4592 = 16'd3959;
parameter WEIGHT_0_4593 = 16'd-3871;
parameter WEIGHT_0_4594 = 16'd428;
parameter WEIGHT_0_4595 = 16'd-5422;
parameter WEIGHT_0_4596 = 16'd13904;
parameter WEIGHT_0_4597 = 16'd-15393;
parameter WEIGHT_0_4598 = 16'd2340;
parameter WEIGHT_0_4599 = 16'd1044;
parameter WEIGHT_0_4600 = 16'd-12112;
parameter WEIGHT_0_4601 = 16'd-439;
parameter WEIGHT_0_4602 = 16'd5727;
parameter WEIGHT_0_4603 = 16'd-1519;
parameter WEIGHT_0_4604 = 16'd1740;
parameter WEIGHT_0_4605 = 16'd-3011;
parameter WEIGHT_0_4606 = 16'd1929;
parameter WEIGHT_0_4607 = 16'd-10563;
parameter WEIGHT_0_4608 = 16'd7584;
parameter WEIGHT_0_4609 = 16'd-1433;
parameter WEIGHT_0_4610 = 16'd-23710;
parameter WEIGHT_0_4611 = 16'd9255;
parameter WEIGHT_0_4612 = 16'd7732;
parameter WEIGHT_0_4613 = 16'd3881;
parameter WEIGHT_0_4614 = 16'd509;
parameter WEIGHT_0_4615 = 16'd-8201;
parameter WEIGHT_0_4616 = 16'd1035;
parameter WEIGHT_0_4617 = 16'd-6528;
parameter WEIGHT_0_4618 = 16'd3433;
parameter WEIGHT_0_4619 = 16'd-6831;
parameter WEIGHT_0_4620 = 16'd-20575;
parameter WEIGHT_0_4621 = 16'd12550;
parameter WEIGHT_0_4622 = 16'd3640;
parameter WEIGHT_0_4623 = 16'd-4568;
parameter WEIGHT_0_4624 = 16'd4225;
parameter WEIGHT_0_4625 = 16'd-8567;
parameter WEIGHT_0_4626 = 16'd2425;
parameter WEIGHT_0_4627 = 16'd-4741;
parameter WEIGHT_0_4628 = 16'd-854;
parameter WEIGHT_0_4629 = 16'd-6385;
parameter WEIGHT_0_4630 = 16'd-17400;
parameter WEIGHT_0_4631 = 16'd1544;
parameter WEIGHT_0_4632 = 16'd427;
parameter WEIGHT_0_4633 = 16'd-6250;
parameter WEIGHT_0_4634 = 16'd13991;
parameter WEIGHT_0_4635 = 16'd-4972;
parameter WEIGHT_0_4636 = 16'd707;
parameter WEIGHT_0_4637 = 16'd174;
parameter WEIGHT_0_4638 = 16'd1071;
parameter WEIGHT_0_4639 = 16'd2476;
parameter WEIGHT_0_4640 = 16'd-7310;
parameter WEIGHT_0_4641 = 16'd-6681;
parameter WEIGHT_0_4642 = 16'd1864;
parameter WEIGHT_0_4643 = 16'd-3356;
parameter WEIGHT_0_4644 = 16'd11519;
parameter WEIGHT_0_4645 = 16'd-4822;
parameter WEIGHT_0_4646 = 16'd-3064;
parameter WEIGHT_0_4647 = 16'd3758;
parameter WEIGHT_0_4648 = 16'd-621;
parameter WEIGHT_0_4649 = 16'd6423;
parameter WEIGHT_0_4650 = 16'd-1505;
parameter WEIGHT_0_4651 = 16'd-19037;
parameter WEIGHT_0_4652 = 16'd2677;
parameter WEIGHT_0_4653 = 16'd-2007;
parameter WEIGHT_0_4654 = 16'd7454;
parameter WEIGHT_0_4655 = 16'd-3625;
parameter WEIGHT_0_4656 = 16'd-3981;
parameter WEIGHT_0_4657 = 16'd4303;
parameter WEIGHT_0_4658 = 16'd-4328;
parameter WEIGHT_0_4659 = 16'd4162;
parameter WEIGHT_0_4660 = 16'd-1199;
parameter WEIGHT_0_4661 = 16'd-15234;
parameter WEIGHT_0_4662 = 16'd-2526;
parameter WEIGHT_0_4663 = 16'd3477;
parameter WEIGHT_0_4664 = 16'd4062;
parameter WEIGHT_0_4665 = 16'd-950;
parameter WEIGHT_0_4666 = 16'd-655;
parameter WEIGHT_0_4667 = 16'd7761;
parameter WEIGHT_0_4668 = 16'd-9912;
parameter WEIGHT_0_4669 = 16'd1964;
parameter WEIGHT_0_4670 = 16'd2430;
parameter WEIGHT_0_4671 = 16'd-15079;
parameter WEIGHT_0_4672 = 16'd751;
parameter WEIGHT_0_4673 = 16'd7551;
parameter WEIGHT_0_4674 = 16'd4177;
parameter WEIGHT_0_4675 = 16'd2040;
parameter WEIGHT_0_4676 = 16'd2903;
parameter WEIGHT_0_4677 = 16'd7413;
parameter WEIGHT_0_4678 = 16'd-8926;
parameter WEIGHT_0_4679 = 16'd-3245;
parameter WEIGHT_0_4680 = 16'd-80;
parameter WEIGHT_0_4681 = 16'd-12208;
parameter WEIGHT_0_4682 = 16'd-761;
parameter WEIGHT_0_4683 = 16'd3263;
parameter WEIGHT_0_4684 = 16'd2950;
parameter WEIGHT_0_4685 = 16'd653;
parameter WEIGHT_0_4686 = 16'd1461;
parameter WEIGHT_0_4687 = 16'd3871;
parameter WEIGHT_0_4688 = 16'd-7992;
parameter WEIGHT_0_4689 = 16'd-3877;
parameter WEIGHT_0_4690 = 16'd2156;
parameter WEIGHT_0_4691 = 16'd-5818;
parameter WEIGHT_0_4692 = 16'd-65;
parameter WEIGHT_0_4693 = 16'd3806;
parameter WEIGHT_0_4694 = 16'd3022;
parameter WEIGHT_0_4695 = 16'd466;
parameter WEIGHT_0_4696 = 16'd313;
parameter WEIGHT_0_4697 = 16'd4826;
parameter WEIGHT_0_4698 = 16'd-8001;
parameter WEIGHT_0_4699 = 16'd-6021;
parameter WEIGHT_0_4700 = 16'd2256;
parameter WEIGHT_0_4701 = 16'd-8254;
parameter WEIGHT_0_4702 = 16'd1951;
parameter WEIGHT_0_4703 = 16'd3693;
parameter WEIGHT_0_4704 = 16'd-425;
parameter WEIGHT_0_4705 = 16'd1272;
parameter WEIGHT_0_4706 = 16'd1830;
parameter WEIGHT_0_4707 = 16'd2593;
parameter WEIGHT_0_4708 = 16'd-11249;
parameter WEIGHT_0_4709 = 16'd-6402;
parameter WEIGHT_0_4710 = 16'd6681;
parameter WEIGHT_0_4711 = 16'd-11033;
parameter WEIGHT_0_4712 = 16'd3106;
parameter WEIGHT_0_4713 = 16'd4059;
parameter WEIGHT_0_4714 = 16'd-6283;
parameter WEIGHT_0_4715 = 16'd1373;
parameter WEIGHT_0_4716 = 16'd507;
parameter WEIGHT_0_4717 = 16'd-1404;
parameter WEIGHT_0_4718 = 16'd-4029;
parameter WEIGHT_0_4719 = 16'd-12225;
parameter WEIGHT_0_4720 = 16'd3357;
parameter WEIGHT_0_4721 = 16'd-5892;
parameter WEIGHT_0_4722 = 16'd9494;
parameter WEIGHT_0_4723 = 16'd4187;
parameter WEIGHT_0_4724 = 16'd-8060;
parameter WEIGHT_0_4725 = 16'd1710;
parameter WEIGHT_0_4726 = 16'd2221;
parameter WEIGHT_0_4727 = 16'd-7834;
parameter WEIGHT_0_4728 = 16'd-5223;
parameter WEIGHT_0_4729 = 16'd-21587;
parameter WEIGHT_0_4730 = 16'd-4900;
parameter WEIGHT_0_4731 = 16'd-8824;
parameter WEIGHT_0_4732 = 16'd18999;
parameter WEIGHT_0_4733 = 16'd-17688;
parameter WEIGHT_0_4734 = 16'd-11730;
parameter WEIGHT_0_4735 = 16'd-8761;
parameter WEIGHT_0_4736 = 16'd-2917;
parameter WEIGHT_0_4737 = 16'd-12975;
parameter WEIGHT_0_4738 = 16'd-10447;
parameter WEIGHT_0_4739 = 16'd-16244;
parameter WEIGHT_0_4740 = 16'd-8186;
parameter WEIGHT_0_4741 = 16'd-6722;
parameter WEIGHT_0_4742 = 16'd14599;
parameter WEIGHT_0_4743 = 16'd-9933;
parameter WEIGHT_0_4744 = 16'd-3929;
parameter WEIGHT_0_4745 = 16'd-13606;
parameter WEIGHT_0_4746 = 16'd-13759;
parameter WEIGHT_0_4747 = 16'd-9677;
parameter WEIGHT_0_4748 = 16'd-11476;
parameter WEIGHT_0_4749 = 16'd-9280;
parameter WEIGHT_0_4750 = 16'd-608;
parameter WEIGHT_0_4751 = 16'd-5262;
parameter WEIGHT_0_4752 = 16'd5950;
parameter WEIGHT_0_4753 = 16'd-5857;
parameter WEIGHT_0_4754 = 16'd-3669;
parameter WEIGHT_0_4755 = 16'd-5009;
parameter WEIGHT_0_4756 = 16'd-2746;
parameter WEIGHT_0_4757 = 16'd-1340;
parameter WEIGHT_0_4758 = 16'd-3877;
parameter WEIGHT_0_4759 = 16'd-4101;
parameter WEIGHT_0_4760 = 16'd-1422;
parameter WEIGHT_0_4761 = 16'd-2077;
parameter WEIGHT_0_4762 = 16'd-1362;
parameter WEIGHT_0_4763 = 16'd453;
parameter WEIGHT_0_4764 = 16'd-2777;
parameter WEIGHT_0_4765 = 16'd2590;
parameter WEIGHT_0_4766 = 16'd2214;
parameter WEIGHT_0_4767 = 16'd1575;
parameter WEIGHT_0_4768 = 16'd-1920;
parameter WEIGHT_0_4769 = 16'd961;
parameter WEIGHT_0_4770 = 16'd784;
parameter WEIGHT_0_4771 = 16'd2756;
parameter WEIGHT_0_4772 = 16'd-3326;
parameter WEIGHT_0_4773 = 16'd5853;
parameter WEIGHT_0_4774 = 16'd1532;
parameter WEIGHT_0_4775 = 16'd-4947;
parameter WEIGHT_0_4776 = 16'd-2632;
parameter WEIGHT_0_4777 = 16'd-5306;
parameter WEIGHT_0_4778 = 16'd-3015;
parameter WEIGHT_0_4779 = 16'd110;
parameter WEIGHT_0_4780 = 16'd-4850;
parameter WEIGHT_0_4781 = 16'd-596;
parameter WEIGHT_0_4782 = 16'd-1035;
parameter WEIGHT_0_4783 = 16'd4089;
parameter WEIGHT_0_4784 = 16'd-3522;
parameter WEIGHT_0_4785 = 16'd-12138;
parameter WEIGHT_0_4786 = 16'd-2258;
parameter WEIGHT_0_4787 = 16'd-4026;
parameter WEIGHT_0_4788 = 16'd-6610;
parameter WEIGHT_0_4789 = 16'd-6672;
parameter WEIGHT_0_4790 = 16'd-6043;
parameter WEIGHT_0_4791 = 16'd-3633;
parameter WEIGHT_0_4792 = 16'd5594;
parameter WEIGHT_0_4793 = 16'd9289;
parameter WEIGHT_0_4794 = 16'd-9377;
parameter WEIGHT_0_4795 = 16'd-163;
parameter WEIGHT_0_4796 = 16'd-13763;
parameter WEIGHT_0_4797 = 16'd-1207;
parameter WEIGHT_0_4798 = 16'd-8832;
parameter WEIGHT_0_4799 = 16'd-6443;
parameter WEIGHT_0_4800 = 16'd-2928;
parameter WEIGHT_0_4801 = 16'd-6974;
parameter WEIGHT_0_4802 = 16'd4778;
parameter WEIGHT_0_4803 = 16'd9364;
parameter WEIGHT_0_4804 = 16'd-4838;
parameter WEIGHT_0_4805 = 16'd-1607;
parameter WEIGHT_0_4806 = 16'd-19195;
parameter WEIGHT_0_4807 = 16'd-121;
parameter WEIGHT_0_4808 = 16'd-9874;
parameter WEIGHT_0_4809 = 16'd-7011;
parameter WEIGHT_0_4810 = 16'd5561;
parameter WEIGHT_0_4811 = 16'd-17035;
parameter WEIGHT_0_4812 = 16'd7556;
parameter WEIGHT_0_4813 = 16'd3596;
parameter WEIGHT_0_4814 = 16'd-5879;
parameter WEIGHT_0_4815 = 16'd4123;
parameter WEIGHT_0_4816 = 16'd-5046;
parameter WEIGHT_0_4817 = 16'd-375;
parameter WEIGHT_0_4818 = 16'd-10268;
parameter WEIGHT_0_4819 = 16'd-5762;
parameter WEIGHT_0_4820 = 16'd4708;
parameter WEIGHT_0_4821 = 16'd-16357;
parameter WEIGHT_0_4822 = 16'd5564;
parameter WEIGHT_0_4823 = 16'd-4940;
parameter WEIGHT_0_4824 = 16'd-1196;
parameter WEIGHT_0_4825 = 16'd4218;
parameter WEIGHT_0_4826 = 16'd-1314;
parameter WEIGHT_0_4827 = 16'd-5347;
parameter WEIGHT_0_4828 = 16'd-7601;
parameter WEIGHT_0_4829 = 16'd-3992;
parameter WEIGHT_0_4830 = 16'd2574;
parameter WEIGHT_0_4831 = 16'd-11430;
parameter WEIGHT_0_4832 = 16'd3585;
parameter WEIGHT_0_4833 = 16'd-4991;
parameter WEIGHT_0_4834 = 16'd4708;
parameter WEIGHT_0_4835 = 16'd-5059;
parameter WEIGHT_0_4836 = 16'd4344;
parameter WEIGHT_0_4837 = 16'd-5481;
parameter WEIGHT_0_4838 = 16'd-943;
parameter WEIGHT_0_4839 = 16'd-1528;
parameter WEIGHT_0_4840 = 16'd4826;
parameter WEIGHT_0_4841 = 16'd-7991;
parameter WEIGHT_0_4842 = 16'd3158;
parameter WEIGHT_0_4843 = 16'd-9655;
parameter WEIGHT_0_4844 = 16'd4121;
parameter WEIGHT_0_4845 = 16'd-9665;
parameter WEIGHT_0_4846 = 16'd6364;
parameter WEIGHT_0_4847 = 16'd-7438;
parameter WEIGHT_0_4848 = 16'd5377;
parameter WEIGHT_0_4849 = 16'd-1274;
parameter WEIGHT_0_4850 = 16'd6450;
parameter WEIGHT_0_4851 = 16'd-6151;
parameter WEIGHT_0_4852 = 16'd829;
parameter WEIGHT_0_4853 = 16'd-11696;
parameter WEIGHT_0_4854 = 16'd1412;
parameter WEIGHT_0_4855 = 16'd-12090;
parameter WEIGHT_0_4856 = 16'd7464;
parameter WEIGHT_0_4857 = 16'd-8127;
parameter WEIGHT_0_4858 = 16'd3837;
parameter WEIGHT_0_4859 = 16'd366;
parameter WEIGHT_0_4860 = 16'd7163;
parameter WEIGHT_0_4861 = 16'd-5215;
parameter WEIGHT_0_4862 = 16'd5037;
parameter WEIGHT_0_4863 = 16'd-14761;
parameter WEIGHT_0_4864 = 16'd639;
parameter WEIGHT_0_4865 = 16'd-10728;
parameter WEIGHT_0_4866 = 16'd9468;
parameter WEIGHT_0_4867 = 16'd-10628;
parameter WEIGHT_0_4868 = 16'd2268;
parameter WEIGHT_0_4869 = 16'd3399;
parameter WEIGHT_0_4870 = 16'd-1549;
parameter WEIGHT_0_4871 = 16'd-3351;
parameter WEIGHT_0_4872 = 16'd6676;
parameter WEIGHT_0_4873 = 16'd-13734;
parameter WEIGHT_0_4874 = 16'd-3910;
parameter WEIGHT_0_4875 = 16'd-10880;
parameter WEIGHT_0_4876 = 16'd10020;
parameter WEIGHT_0_4877 = 16'd-8324;
parameter WEIGHT_0_4878 = 16'd6415;
parameter WEIGHT_0_4879 = 16'd522;
parameter WEIGHT_0_4880 = 16'd-7440;
parameter WEIGHT_0_4881 = 16'd272;
parameter WEIGHT_0_4882 = 16'd7955;
parameter WEIGHT_0_4883 = 16'd-9529;
parameter WEIGHT_0_4884 = 16'd2554;
parameter WEIGHT_0_4885 = 16'd-12674;
parameter WEIGHT_0_4886 = 16'd3834;
parameter WEIGHT_0_4887 = 16'd-4090;
parameter WEIGHT_0_4888 = 16'd8406;
parameter WEIGHT_0_4889 = 16'd-2095;
parameter WEIGHT_0_4890 = 16'd-19335;
parameter WEIGHT_0_4891 = 16'd8628;
parameter WEIGHT_0_4892 = 16'd4950;
parameter WEIGHT_0_4893 = 16'd-9213;
parameter WEIGHT_0_4894 = 16'd4164;
parameter WEIGHT_0_4895 = 16'd-9602;
parameter WEIGHT_0_4896 = 16'd1057;
parameter WEIGHT_0_4897 = 16'd-62;
parameter WEIGHT_0_4898 = 16'd2757;
parameter WEIGHT_0_4899 = 16'd-3466;
parameter WEIGHT_0_4900 = 16'd-18959;
parameter WEIGHT_0_4901 = 16'd10191;
parameter WEIGHT_0_4902 = 16'd1924;
parameter WEIGHT_0_4903 = 16'd-10066;
parameter WEIGHT_0_4904 = 16'd10610;
parameter WEIGHT_0_4905 = 16'd-8891;
parameter WEIGHT_0_4906 = 16'd-107;
parameter WEIGHT_0_4907 = 16'd186;
parameter WEIGHT_0_4908 = 16'd-2087;
parameter WEIGHT_0_4909 = 16'd-2937;
parameter WEIGHT_0_4910 = 16'd-10068;
parameter WEIGHT_0_4911 = 16'd1346;
parameter WEIGHT_0_4912 = 16'd-541;
parameter WEIGHT_0_4913 = 16'd-6353;
parameter WEIGHT_0_4914 = 16'd9475;
parameter WEIGHT_0_4915 = 16'd-4771;
parameter WEIGHT_0_4916 = 16'd-1524;
parameter WEIGHT_0_4917 = 16'd2301;
parameter WEIGHT_0_4918 = 16'd-3918;
parameter WEIGHT_0_4919 = 16'd2627;
parameter WEIGHT_0_4920 = 16'd-4850;
parameter WEIGHT_0_4921 = 16'd-10680;
parameter WEIGHT_0_4922 = 16'd2593;
parameter WEIGHT_0_4923 = 16'd-48;
parameter WEIGHT_0_4924 = 16'd7800;
parameter WEIGHT_0_4925 = 16'd-1477;
parameter WEIGHT_0_4926 = 16'd-3958;
parameter WEIGHT_0_4927 = 16'd435;
parameter WEIGHT_0_4928 = 16'd-2265;
parameter WEIGHT_0_4929 = 16'd559;
parameter WEIGHT_0_4930 = 16'd792;
parameter WEIGHT_0_4931 = 16'd-11976;
parameter WEIGHT_0_4932 = 16'd1335;
parameter WEIGHT_0_4933 = 16'd3855;
parameter WEIGHT_0_4934 = 16'd5446;
parameter WEIGHT_0_4935 = 16'd2809;
parameter WEIGHT_0_4936 = 16'd721;
parameter WEIGHT_0_4937 = 16'd2558;
parameter WEIGHT_0_4938 = 16'd-3197;
parameter WEIGHT_0_4939 = 16'd-1112;
parameter WEIGHT_0_4940 = 16'd-1733;
parameter WEIGHT_0_4941 = 16'd-12033;
parameter WEIGHT_0_4942 = 16'd-896;
parameter WEIGHT_0_4943 = 16'd1941;
parameter WEIGHT_0_4944 = 16'd1331;
parameter WEIGHT_0_4945 = 16'd1026;
parameter WEIGHT_0_4946 = 16'd1953;
parameter WEIGHT_0_4947 = 16'd-22;
parameter WEIGHT_0_4948 = 16'd-5236;
parameter WEIGHT_0_4949 = 16'd-2508;
parameter WEIGHT_0_4950 = 16'd2334;
parameter WEIGHT_0_4951 = 16'd-8685;
parameter WEIGHT_0_4952 = 16'd-716;
parameter WEIGHT_0_4953 = 16'd5626;
parameter WEIGHT_0_4954 = 16'd-775;
parameter WEIGHT_0_4955 = 16'd1317;
parameter WEIGHT_0_4956 = 16'd1662;
parameter WEIGHT_0_4957 = 16'd2108;
parameter WEIGHT_0_4958 = 16'd-6355;
parameter WEIGHT_0_4959 = 16'd-2901;
parameter WEIGHT_0_4960 = 16'd3362;
parameter WEIGHT_0_4961 = 16'd-4821;
parameter WEIGHT_0_4962 = 16'd518;
parameter WEIGHT_0_4963 = 16'd811;
parameter WEIGHT_0_4964 = 16'd-2820;
parameter WEIGHT_0_4965 = 16'd-72;
parameter WEIGHT_0_4966 = 16'd-63;
parameter WEIGHT_0_4967 = 16'd95;
parameter WEIGHT_0_4968 = 16'd-5182;
parameter WEIGHT_0_4969 = 16'd-6157;
parameter WEIGHT_0_4970 = 16'd2761;
parameter WEIGHT_0_4971 = 16'd-3106;
parameter WEIGHT_0_4972 = 16'd1953;
parameter WEIGHT_0_4973 = 16'd5100;
parameter WEIGHT_0_4974 = 16'd-21;
parameter WEIGHT_0_4975 = 16'd-460;
parameter WEIGHT_0_4976 = 16'd284;
parameter WEIGHT_0_4977 = 16'd-1366;
parameter WEIGHT_0_4978 = 16'd-6553;
parameter WEIGHT_0_4979 = 16'd-6938;
parameter WEIGHT_0_4980 = 16'd4776;
parameter WEIGHT_0_4981 = 16'd-5812;
parameter WEIGHT_0_4982 = 16'd3325;
parameter WEIGHT_0_4983 = 16'd6296;
parameter WEIGHT_0_4984 = 16'd-3784;
parameter WEIGHT_0_4985 = 16'd-1616;
parameter WEIGHT_0_4986 = 16'd-1975;
parameter WEIGHT_0_4987 = 16'd-3006;
parameter WEIGHT_0_4988 = 16'd-5793;
parameter WEIGHT_0_4989 = 16'd-10480;
parameter WEIGHT_0_4990 = 16'd370;
parameter WEIGHT_0_4991 = 16'd-7127;
parameter WEIGHT_0_4992 = 16'd4258;
parameter WEIGHT_0_4993 = 16'd5582;
parameter WEIGHT_0_4994 = 16'd-7856;
parameter WEIGHT_0_4995 = 16'd3478;
parameter WEIGHT_0_4996 = 16'd-1474;
parameter WEIGHT_0_4997 = 16'd-7689;
parameter WEIGHT_0_4998 = 16'd-3116;
parameter WEIGHT_0_4999 = 16'd-15436;
parameter WEIGHT_0_5000 = 16'd-1632;
parameter WEIGHT_0_5001 = 16'd-3430;
parameter WEIGHT_0_5002 = 16'd11990;
parameter WEIGHT_0_5003 = 16'd-3845;
parameter WEIGHT_0_5004 = 16'd-9179;
parameter WEIGHT_0_5005 = 16'd4332;
parameter WEIGHT_0_5006 = 16'd-739;
parameter WEIGHT_0_5007 = 16'd-1174;
parameter WEIGHT_0_5008 = 16'd907;
parameter WEIGHT_0_5009 = 16'd-20837;
parameter WEIGHT_0_5010 = 16'd-7319;
parameter WEIGHT_0_5011 = 16'd-11283;
parameter WEIGHT_0_5012 = 16'd18809;
parameter WEIGHT_0_5013 = 16'd-14545;
parameter WEIGHT_0_5014 = 16'd-11004;
parameter WEIGHT_0_5015 = 16'd-10322;
parameter WEIGHT_0_5016 = 16'd-5811;
parameter WEIGHT_0_5017 = 16'd271;
parameter WEIGHT_0_5018 = 16'd-21038;
parameter WEIGHT_0_5019 = 16'd-11378;
parameter WEIGHT_0_5020 = 16'd-5250;
parameter WEIGHT_0_5021 = 16'd-6473;
parameter WEIGHT_0_5022 = 16'd10354;
parameter WEIGHT_0_5023 = 16'd-8850;
parameter WEIGHT_0_5024 = 16'd-8404;
parameter WEIGHT_0_5025 = 16'd-12256;
parameter WEIGHT_0_5026 = 16'd-11278;
parameter WEIGHT_0_5027 = 16'd-2309;
parameter WEIGHT_0_5028 = 16'd-9191;
parameter WEIGHT_0_5029 = 16'd-8683;
parameter WEIGHT_0_5030 = 16'd-1501;
parameter WEIGHT_0_5031 = 16'd-3114;
parameter WEIGHT_0_5032 = 16'd7528;
parameter WEIGHT_0_5033 = 16'd-3637;
parameter WEIGHT_0_5034 = 16'd-5386;
parameter WEIGHT_0_5035 = 16'd-6606;
parameter WEIGHT_0_5036 = 16'd-9578;
parameter WEIGHT_0_5037 = 16'd-3720;
parameter WEIGHT_0_5038 = 16'd-6926;
parameter WEIGHT_0_5039 = 16'd-4962;
parameter WEIGHT_0_5040 = 16'd-163;
parameter WEIGHT_0_5041 = 16'd-2730;
parameter WEIGHT_0_5042 = 16'd-5980;
parameter WEIGHT_0_5043 = 16'd-2783;
parameter WEIGHT_0_5044 = 16'd-4433;
parameter WEIGHT_0_5045 = 16'd-1759;
parameter WEIGHT_0_5046 = 16'd-4072;
parameter WEIGHT_0_5047 = 16'd3588;
parameter WEIGHT_0_5048 = 16'd-2607;
parameter WEIGHT_0_5049 = 16'd446;
parameter WEIGHT_0_5050 = 16'd-817;
parameter WEIGHT_0_5051 = 16'd4760;
parameter WEIGHT_0_5052 = 16'd-4337;
parameter WEIGHT_0_5053 = 16'd1782;
parameter WEIGHT_0_5054 = 16'd-2081;
parameter WEIGHT_0_5055 = 16'd-5014;
parameter WEIGHT_0_5056 = 16'd1676;
parameter WEIGHT_0_5057 = 16'd-510;
parameter WEIGHT_0_5058 = 16'd-3508;
parameter WEIGHT_0_5059 = 16'd-2514;
parameter WEIGHT_0_5060 = 16'd-8011;
parameter WEIGHT_0_5061 = 16'd-783;
parameter WEIGHT_0_5062 = 16'd-4721;
parameter WEIGHT_0_5063 = 16'd5020;
parameter WEIGHT_0_5064 = 16'd-5714;
parameter WEIGHT_0_5065 = 16'd-7668;
parameter WEIGHT_0_5066 = 16'd-1435;
parameter WEIGHT_0_5067 = 16'd2792;
parameter WEIGHT_0_5068 = 16'd-6100;
parameter WEIGHT_0_5069 = 16'd-9659;
parameter WEIGHT_0_5070 = 16'd-12349;
parameter WEIGHT_0_5071 = 16'd-1782;
parameter WEIGHT_0_5072 = 16'd-115;
parameter WEIGHT_0_5073 = 16'd11865;
parameter WEIGHT_0_5074 = 16'd-10677;
parameter WEIGHT_0_5075 = 16'd1502;
parameter WEIGHT_0_5076 = 16'd-9554;
parameter WEIGHT_0_5077 = 16'd-197;
parameter WEIGHT_0_5078 = 16'd-18451;
parameter WEIGHT_0_5079 = 16'd-11812;
parameter WEIGHT_0_5080 = 16'd-3980;
parameter WEIGHT_0_5081 = 16'd-13978;
parameter WEIGHT_0_5082 = 16'd8366;
parameter WEIGHT_0_5083 = 16'd6890;
parameter WEIGHT_0_5084 = 16'd-8029;
parameter WEIGHT_0_5085 = 16'd2438;
parameter WEIGHT_0_5086 = 16'd-16194;
parameter WEIGHT_0_5087 = 16'd-4238;
parameter WEIGHT_0_5088 = 16'd-10397;
parameter WEIGHT_0_5089 = 16'd-9394;
parameter WEIGHT_0_5090 = 16'd-1051;
parameter WEIGHT_0_5091 = 16'd-21508;
parameter WEIGHT_0_5092 = 16'd7237;
parameter WEIGHT_0_5093 = 16'd6990;
parameter WEIGHT_0_5094 = 16'd-7205;
parameter WEIGHT_0_5095 = 16'd7502;
parameter WEIGHT_0_5096 = 16'd-11160;
parameter WEIGHT_0_5097 = 16'd-6132;
parameter WEIGHT_0_5098 = 16'd-4600;
parameter WEIGHT_0_5099 = 16'd-7015;
parameter WEIGHT_0_5100 = 16'd1618;
parameter WEIGHT_0_5101 = 16'd-18993;
parameter WEIGHT_0_5102 = 16'd3821;
parameter WEIGHT_0_5103 = 16'd3447;
parameter WEIGHT_0_5104 = 16'd-4997;
parameter WEIGHT_0_5105 = 16'd7185;
parameter WEIGHT_0_5106 = 16'd-3006;
parameter WEIGHT_0_5107 = 16'd-10522;
parameter WEIGHT_0_5108 = 16'd-1153;
parameter WEIGHT_0_5109 = 16'd-909;
parameter WEIGHT_0_5110 = 16'd3888;
parameter WEIGHT_0_5111 = 16'd-12757;
parameter WEIGHT_0_5112 = 16'd5697;
parameter WEIGHT_0_5113 = 16'd-3777;
parameter WEIGHT_0_5114 = 16'd-1357;
parameter WEIGHT_0_5115 = 16'd4890;
parameter WEIGHT_0_5116 = 16'd63;
parameter WEIGHT_0_5117 = 16'd-9592;
parameter WEIGHT_0_5118 = 16'd-594;
parameter WEIGHT_0_5119 = 16'd-4566;
parameter WEIGHT_0_5120 = 16'd4158;
parameter WEIGHT_0_5121 = 16'd-5180;
parameter WEIGHT_0_5122 = 16'd1369;
parameter WEIGHT_0_5123 = 16'd-5822;
parameter WEIGHT_0_5124 = 16'd-2457;
parameter WEIGHT_0_5125 = 16'd-4033;
parameter WEIGHT_0_5126 = 16'd1740;
parameter WEIGHT_0_5127 = 16'd-10576;
parameter WEIGHT_0_5128 = 16'd4529;
parameter WEIGHT_0_5129 = 16'd108;
parameter WEIGHT_0_5130 = 16'd5228;
parameter WEIGHT_0_5131 = 16'd337;
parameter WEIGHT_0_5132 = 16'd4200;
parameter WEIGHT_0_5133 = 16'd-10045;
parameter WEIGHT_0_5134 = 16'd-2080;
parameter WEIGHT_0_5135 = 16'd-6401;
parameter WEIGHT_0_5136 = 16'd4546;
parameter WEIGHT_0_5137 = 16'd-11161;
parameter WEIGHT_0_5138 = 16'd7724;
parameter WEIGHT_0_5139 = 16'd1934;
parameter WEIGHT_0_5140 = 16'd7587;
parameter WEIGHT_0_5141 = 16'd-3731;
parameter WEIGHT_0_5142 = 16'd3618;
parameter WEIGHT_0_5143 = 16'd-15102;
parameter WEIGHT_0_5144 = 16'd-8316;
parameter WEIGHT_0_5145 = 16'd-8186;
parameter WEIGHT_0_5146 = 16'd10511;
parameter WEIGHT_0_5147 = 16'd-13038;
parameter WEIGHT_0_5148 = 16'd3536;
parameter WEIGHT_0_5149 = 16'd192;
parameter WEIGHT_0_5150 = 16'd1118;
parameter WEIGHT_0_5151 = 16'd-4254;
parameter WEIGHT_0_5152 = 16'd3954;
parameter WEIGHT_0_5153 = 16'd-13207;
parameter WEIGHT_0_5154 = 16'd-3973;
parameter WEIGHT_0_5155 = 16'd-6897;
parameter WEIGHT_0_5156 = 16'd10030;
parameter WEIGHT_0_5157 = 16'd-8468;
parameter WEIGHT_0_5158 = 16'd5740;
parameter WEIGHT_0_5159 = 16'd-2305;
parameter WEIGHT_0_5160 = 16'd-9602;
parameter WEIGHT_0_5161 = 16'd1524;
parameter WEIGHT_0_5162 = 16'd6522;
parameter WEIGHT_0_5163 = 16'd-12837;
parameter WEIGHT_0_5164 = 16'd-637;
parameter WEIGHT_0_5165 = 16'd-7707;
parameter WEIGHT_0_5166 = 16'd7976;
parameter WEIGHT_0_5167 = 16'd-3467;
parameter WEIGHT_0_5168 = 16'd1942;
parameter WEIGHT_0_5169 = 16'd-7489;
parameter WEIGHT_0_5170 = 16'd-17186;
parameter WEIGHT_0_5171 = 16'd8164;
parameter WEIGHT_0_5172 = 16'd4777;
parameter WEIGHT_0_5173 = 16'd-13370;
parameter WEIGHT_0_5174 = 16'd2996;
parameter WEIGHT_0_5175 = 16'd-4065;
parameter WEIGHT_0_5176 = 16'd4515;
parameter WEIGHT_0_5177 = 16'd341;
parameter WEIGHT_0_5178 = 16'd-2582;
parameter WEIGHT_0_5179 = 16'd-5583;
parameter WEIGHT_0_5180 = 16'd-15022;
parameter WEIGHT_0_5181 = 16'd8204;
parameter WEIGHT_0_5182 = 16'd3281;
parameter WEIGHT_0_5183 = 16'd-9028;
parameter WEIGHT_0_5184 = 16'd7876;
parameter WEIGHT_0_5185 = 16'd-1377;
parameter WEIGHT_0_5186 = 16'd651;
parameter WEIGHT_0_5187 = 16'd2387;
parameter WEIGHT_0_5188 = 16'd-3955;
parameter WEIGHT_0_5189 = 16'd-828;
parameter WEIGHT_0_5190 = 16'd-3918;
parameter WEIGHT_0_5191 = 16'd-1838;
parameter WEIGHT_0_5192 = 16'd2984;
parameter WEIGHT_0_5193 = 16'd-1969;
parameter WEIGHT_0_5194 = 16'd7186;
parameter WEIGHT_0_5195 = 16'd879;
parameter WEIGHT_0_5196 = 16'd2207;
parameter WEIGHT_0_5197 = 16'd234;
parameter WEIGHT_0_5198 = 16'd-1616;
parameter WEIGHT_0_5199 = 16'd2256;
parameter WEIGHT_0_5200 = 16'd-3462;
parameter WEIGHT_0_5201 = 16'd-9271;
parameter WEIGHT_0_5202 = 16'd1205;
parameter WEIGHT_0_5203 = 16'd4522;
parameter WEIGHT_0_5204 = 16'd6760;
parameter WEIGHT_0_5205 = 16'd1226;
parameter WEIGHT_0_5206 = 16'd3192;
parameter WEIGHT_0_5207 = 16'd-3647;
parameter WEIGHT_0_5208 = 16'd-1578;
parameter WEIGHT_0_5209 = 16'd-815;
parameter WEIGHT_0_5210 = 16'd-970;
parameter WEIGHT_0_5211 = 16'd-6811;
parameter WEIGHT_0_5212 = 16'd2711;
parameter WEIGHT_0_5213 = 16'd5367;
parameter WEIGHT_0_5214 = 16'd-3426;
parameter WEIGHT_0_5215 = 16'd2238;
parameter WEIGHT_0_5216 = 16'd4799;
parameter WEIGHT_0_5217 = 16'd-3647;
parameter WEIGHT_0_5218 = 16'd-3354;
parameter WEIGHT_0_5219 = 16'd224;
parameter WEIGHT_0_5220 = 16'd-1594;
parameter WEIGHT_0_5221 = 16'd-6624;
parameter WEIGHT_0_5222 = 16'd3796;
parameter WEIGHT_0_5223 = 16'd5751;
parameter WEIGHT_0_5224 = 16'd-1921;
parameter WEIGHT_0_5225 = 16'd770;
parameter WEIGHT_0_5226 = 16'd3608;
parameter WEIGHT_0_5227 = 16'd-1643;
parameter WEIGHT_0_5228 = 16'd-2590;
parameter WEIGHT_0_5229 = 16'd-2912;
parameter WEIGHT_0_5230 = 16'd-2928;
parameter WEIGHT_0_5231 = 16'd-1508;
parameter WEIGHT_0_5232 = 16'd-23;
parameter WEIGHT_0_5233 = 16'd3777;
parameter WEIGHT_0_5234 = 16'd-2465;
parameter WEIGHT_0_5235 = 16'd-290;
parameter WEIGHT_0_5236 = 16'd3119;
parameter WEIGHT_0_5237 = 16'd-4562;
parameter WEIGHT_0_5238 = 16'd-4116;
parameter WEIGHT_0_5239 = 16'd-4619;
parameter WEIGHT_0_5240 = 16'd-1625;
parameter WEIGHT_0_5241 = 16'd-2653;
parameter WEIGHT_0_5242 = 16'd-826;
parameter WEIGHT_0_5243 = 16'd5868;
parameter WEIGHT_0_5244 = 16'd-2067;
parameter WEIGHT_0_5245 = 16'd2627;
parameter WEIGHT_0_5246 = 16'd-1741;
parameter WEIGHT_0_5247 = 16'd-1770;
parameter WEIGHT_0_5248 = 16'd-2653;
parameter WEIGHT_0_5249 = 16'd-1642;
parameter WEIGHT_0_5250 = 16'd-1090;
parameter WEIGHT_0_5251 = 16'd187;
parameter WEIGHT_0_5252 = 16'd2883;
parameter WEIGHT_0_5253 = 16'd7948;
parameter WEIGHT_0_5254 = 16'd-5750;
parameter WEIGHT_0_5255 = 16'd2732;
parameter WEIGHT_0_5256 = 16'd2098;
parameter WEIGHT_0_5257 = 16'd-4778;
parameter WEIGHT_0_5258 = 16'd-1671;
parameter WEIGHT_0_5259 = 16'd-6290;
parameter WEIGHT_0_5260 = 16'd1210;
parameter WEIGHT_0_5261 = 16'd-3557;
parameter WEIGHT_0_5262 = 16'd3413;
parameter WEIGHT_0_5263 = 16'd4852;
parameter WEIGHT_0_5264 = 16'd-9521;
parameter WEIGHT_0_5265 = 16'd2219;
parameter WEIGHT_0_5266 = 16'd-3450;
parameter WEIGHT_0_5267 = 16'd-9269;
parameter WEIGHT_0_5268 = 16'd-2311;
parameter WEIGHT_0_5269 = 16'd-10364;
parameter WEIGHT_0_5270 = 16'd-479;
parameter WEIGHT_0_5271 = 16'd-6827;
parameter WEIGHT_0_5272 = 16'd9459;
parameter WEIGHT_0_5273 = 16'd2732;
parameter WEIGHT_0_5274 = 16'd-7916;
parameter WEIGHT_0_5275 = 16'd1762;
parameter WEIGHT_0_5276 = 16'd1078;
parameter WEIGHT_0_5277 = 16'd-13532;
parameter WEIGHT_0_5278 = 16'd1839;
parameter WEIGHT_0_5279 = 16'd-13249;
parameter WEIGHT_0_5280 = 16'd-3750;
parameter WEIGHT_0_5281 = 16'd-608;
parameter WEIGHT_0_5282 = 16'd13746;
parameter WEIGHT_0_5283 = 16'd-10578;
parameter WEIGHT_0_5284 = 16'd-11148;
parameter WEIGHT_0_5285 = 16'd2757;
parameter WEIGHT_0_5286 = 16'd-3630;
parameter WEIGHT_0_5287 = 16'd-6172;
parameter WEIGHT_0_5288 = 16'd-4726;
parameter WEIGHT_0_5289 = 16'd-15561;
parameter WEIGHT_0_5290 = 16'd-6766;
parameter WEIGHT_0_5291 = 16'd-5401;
parameter WEIGHT_0_5292 = 16'd15397;
parameter WEIGHT_0_5293 = 16'd-18138;
parameter WEIGHT_0_5294 = 16'd-14779;
parameter WEIGHT_0_5295 = 16'd-7041;
parameter WEIGHT_0_5296 = 16'd-2050;
parameter WEIGHT_0_5297 = 16'd-4679;
parameter WEIGHT_0_5298 = 16'd-16686;
parameter WEIGHT_0_5299 = 16'd-11984;
parameter WEIGHT_0_5300 = 16'd-5047;
parameter WEIGHT_0_5301 = 16'd-1294;
parameter WEIGHT_0_5302 = 16'd8397;
parameter WEIGHT_0_5303 = 16'd-11210;
parameter WEIGHT_0_5304 = 16'd-2100;
parameter WEIGHT_0_5305 = 16'd-8765;
parameter WEIGHT_0_5306 = 16'd-4110;
parameter WEIGHT_0_5307 = 16'd-279;
parameter WEIGHT_0_5308 = 16'd-6980;
parameter WEIGHT_0_5309 = 16'd-7079;
parameter WEIGHT_0_5310 = 16'd-3798;
parameter WEIGHT_0_5311 = 16'd3470;
parameter WEIGHT_0_5312 = 16'd4895;
parameter WEIGHT_0_5313 = 16'd-6720;
parameter WEIGHT_0_5314 = 16'd-4601;
parameter WEIGHT_0_5315 = 16'd-2637;
parameter WEIGHT_0_5316 = 16'd-7765;
parameter WEIGHT_0_5317 = 16'd-2773;
parameter WEIGHT_0_5318 = 16'd-3368;
parameter WEIGHT_0_5319 = 16'd-5543;
parameter WEIGHT_0_5320 = 16'd804;
parameter WEIGHT_0_5321 = 16'd2275;
parameter WEIGHT_0_5322 = 16'd-2135;
parameter WEIGHT_0_5323 = 16'd-957;
parameter WEIGHT_0_5324 = 16'd135;
parameter WEIGHT_0_5325 = 16'd1133;
parameter WEIGHT_0_5326 = 16'd-1518;
parameter WEIGHT_0_5327 = 16'd-106;
parameter WEIGHT_0_5328 = 16'd-2660;
parameter WEIGHT_0_5329 = 16'd329;
parameter WEIGHT_0_5330 = 16'd-552;
parameter WEIGHT_0_5331 = 16'd624;
parameter WEIGHT_0_5332 = 16'd-5398;
parameter WEIGHT_0_5333 = 16'd1180;
parameter WEIGHT_0_5334 = 16'd-4735;
parameter WEIGHT_0_5335 = 16'd-5550;
parameter WEIGHT_0_5336 = 16'd-2216;
parameter WEIGHT_0_5337 = 16'd2378;
parameter WEIGHT_0_5338 = 16'd-6435;
parameter WEIGHT_0_5339 = 16'd-5767;
parameter WEIGHT_0_5340 = 16'd-3623;
parameter WEIGHT_0_5341 = 16'd-3849;
parameter WEIGHT_0_5342 = 16'd-6492;
parameter WEIGHT_0_5343 = 16'd17;
parameter WEIGHT_0_5344 = 16'd-4329;
parameter WEIGHT_0_5345 = 16'd604;
parameter WEIGHT_0_5346 = 16'd-590;
parameter WEIGHT_0_5347 = 16'd4918;
parameter WEIGHT_0_5348 = 16'd-6467;
parameter WEIGHT_0_5349 = 16'd-10710;
parameter WEIGHT_0_5350 = 16'd-10232;
parameter WEIGHT_0_5351 = 16'd-8167;
parameter WEIGHT_0_5352 = 16'd-4305;
parameter WEIGHT_0_5353 = 16'd12737;
parameter WEIGHT_0_5354 = 16'd-5879;
parameter WEIGHT_0_5355 = 16'd-2147;
parameter WEIGHT_0_5356 = 16'd-12174;
parameter WEIGHT_0_5357 = 16'd-1296;
parameter WEIGHT_0_5358 = 16'd-16533;
parameter WEIGHT_0_5359 = 16'd-11192;
parameter WEIGHT_0_5360 = 16'd-3927;
parameter WEIGHT_0_5361 = 16'd-15094;
parameter WEIGHT_0_5362 = 16'd4724;
parameter WEIGHT_0_5363 = 16'd8811;
parameter WEIGHT_0_5364 = 16'd-8197;
parameter WEIGHT_0_5365 = 16'd3229;
parameter WEIGHT_0_5366 = 16'd-13867;
parameter WEIGHT_0_5367 = 16'd-4044;
parameter WEIGHT_0_5368 = 16'd-8465;
parameter WEIGHT_0_5369 = 16'd-12414;
parameter WEIGHT_0_5370 = 16'd-271;
parameter WEIGHT_0_5371 = 16'd-21327;
parameter WEIGHT_0_5372 = 16'd3500;
parameter WEIGHT_0_5373 = 16'd7821;
parameter WEIGHT_0_5374 = 16'd-5733;
parameter WEIGHT_0_5375 = 16'd4374;
parameter WEIGHT_0_5376 = 16'd-10847;
parameter WEIGHT_0_5377 = 16'd-6328;
parameter WEIGHT_0_5378 = 16'd-2291;
parameter WEIGHT_0_5379 = 16'd-6198;
parameter WEIGHT_0_5380 = 16'd752;
parameter WEIGHT_0_5381 = 16'd-11612;
parameter WEIGHT_0_5382 = 16'd5710;
parameter WEIGHT_0_5383 = 16'd5299;
parameter WEIGHT_0_5384 = 16'd-7678;
parameter WEIGHT_0_5385 = 16'd8553;
parameter WEIGHT_0_5386 = 16'd-7357;
parameter WEIGHT_0_5387 = 16'd-13366;
parameter WEIGHT_0_5388 = 16'd-180;
parameter WEIGHT_0_5389 = 16'd-8280;
parameter WEIGHT_0_5390 = 16'd2641;
parameter WEIGHT_0_5391 = 16'd-6462;
parameter WEIGHT_0_5392 = 16'd4064;
parameter WEIGHT_0_5393 = 16'd3689;
parameter WEIGHT_0_5394 = 16'd-8648;
parameter WEIGHT_0_5395 = 16'd6318;
parameter WEIGHT_0_5396 = 16'd-3229;
parameter WEIGHT_0_5397 = 16'd-13385;
parameter WEIGHT_0_5398 = 16'd506;
parameter WEIGHT_0_5399 = 16'd-1995;
parameter WEIGHT_0_5400 = 16'd1499;
parameter WEIGHT_0_5401 = 16'd-860;
parameter WEIGHT_0_5402 = 16'd7181;
parameter WEIGHT_0_5403 = 16'd-3032;
parameter WEIGHT_0_5404 = 16'd-9094;
parameter WEIGHT_0_5405 = 16'd5391;
parameter WEIGHT_0_5406 = 16'd2130;
parameter WEIGHT_0_5407 = 16'd-10424;
parameter WEIGHT_0_5408 = 16'd-1074;
parameter WEIGHT_0_5409 = 16'd-6995;
parameter WEIGHT_0_5410 = 16'd5726;
parameter WEIGHT_0_5411 = 16'd215;
parameter WEIGHT_0_5412 = 16'd3194;
parameter WEIGHT_0_5413 = 16'd-1650;
parameter WEIGHT_0_5414 = 16'd-13496;
parameter WEIGHT_0_5415 = 16'd1880;
parameter WEIGHT_0_5416 = 16'd5105;
parameter WEIGHT_0_5417 = 16'd-8897;
parameter WEIGHT_0_5418 = 16'd3185;
parameter WEIGHT_0_5419 = 16'd-10131;
parameter WEIGHT_0_5420 = 16'd6868;
parameter WEIGHT_0_5421 = 16'd-2856;
parameter WEIGHT_0_5422 = 16'd3869;
parameter WEIGHT_0_5423 = 16'd-7648;
parameter WEIGHT_0_5424 = 16'd-13965;
parameter WEIGHT_0_5425 = 16'd-3080;
parameter WEIGHT_0_5426 = 16'd6317;
parameter WEIGHT_0_5427 = 16'd-7563;
parameter WEIGHT_0_5428 = 16'd2658;
parameter WEIGHT_0_5429 = 16'd-7448;
parameter WEIGHT_0_5430 = 16'd4032;
parameter WEIGHT_0_5431 = 16'd-21;
parameter WEIGHT_0_5432 = 16'd7468;
parameter WEIGHT_0_5433 = 16'd-7741;
parameter WEIGHT_0_5434 = 16'd-9941;
parameter WEIGHT_0_5435 = 16'd-2244;
parameter WEIGHT_0_5436 = 16'd10210;
parameter WEIGHT_0_5437 = 16'd-7065;
parameter WEIGHT_0_5438 = 16'd-2494;
parameter WEIGHT_0_5439 = 16'd-7619;
parameter WEIGHT_0_5440 = 16'd-464;
parameter WEIGHT_0_5441 = 16'd276;
parameter WEIGHT_0_5442 = 16'd5033;
parameter WEIGHT_0_5443 = 16'd-9418;
parameter WEIGHT_0_5444 = 16'd-6960;
parameter WEIGHT_0_5445 = 16'd1970;
parameter WEIGHT_0_5446 = 16'd12291;
parameter WEIGHT_0_5447 = 16'd-2975;
parameter WEIGHT_0_5448 = 16'd-1676;
parameter WEIGHT_0_5449 = 16'd-10459;
parameter WEIGHT_0_5450 = 16'd-5860;
parameter WEIGHT_0_5451 = 16'd6681;
parameter WEIGHT_0_5452 = 16'd7259;
parameter WEIGHT_0_5453 = 16'd-7791;
parameter WEIGHT_0_5454 = 16'd-1788;
parameter WEIGHT_0_5455 = 16'd-912;
parameter WEIGHT_0_5456 = 16'd2945;
parameter WEIGHT_0_5457 = 16'd1672;
parameter WEIGHT_0_5458 = 16'd-3814;
parameter WEIGHT_0_5459 = 16'd-6106;
parameter WEIGHT_0_5460 = 16'd-3579;
parameter WEIGHT_0_5461 = 16'd1530;
parameter WEIGHT_0_5462 = 16'd1641;
parameter WEIGHT_0_5463 = 16'd-1723;
parameter WEIGHT_0_5464 = 16'd604;
parameter WEIGHT_0_5465 = 16'd186;
parameter WEIGHT_0_5466 = 16'd5031;
parameter WEIGHT_0_5467 = 16'd1084;
parameter WEIGHT_0_5468 = 16'd-6210;
parameter WEIGHT_0_5469 = 16'd-1193;
parameter WEIGHT_0_5470 = 16'd-2322;
parameter WEIGHT_0_5471 = 16'd-1302;
parameter WEIGHT_0_5472 = 16'd1093;
parameter WEIGHT_0_5473 = 16'd1005;
parameter WEIGHT_0_5474 = 16'd1336;
parameter WEIGHT_0_5475 = 16'd1457;
parameter WEIGHT_0_5476 = 16'd3152;
parameter WEIGHT_0_5477 = 16'd-2055;
parameter WEIGHT_0_5478 = 16'd-4283;
parameter WEIGHT_0_5479 = 16'd-3199;
parameter WEIGHT_0_5480 = 16'd-910;
parameter WEIGHT_0_5481 = 16'd161;
parameter WEIGHT_0_5482 = 16'd3307;
parameter WEIGHT_0_5483 = 16'd2368;
parameter WEIGHT_0_5484 = 16'd-1660;
parameter WEIGHT_0_5485 = 16'd-1164;
parameter WEIGHT_0_5486 = 16'd6454;
parameter WEIGHT_0_5487 = 16'd-3372;
parameter WEIGHT_0_5488 = 16'd-1125;
parameter WEIGHT_0_5489 = 16'd-2696;
parameter WEIGHT_0_5490 = 16'd2104;
parameter WEIGHT_0_5491 = 16'd-2369;
parameter WEIGHT_0_5492 = 16'd2096;
parameter WEIGHT_0_5493 = 16'd7899;
parameter WEIGHT_0_5494 = 16'd-2501;
parameter WEIGHT_0_5495 = 16'd1920;
parameter WEIGHT_0_5496 = 16'd5777;
parameter WEIGHT_0_5497 = 16'd-4758;
parameter WEIGHT_0_5498 = 16'd-960;
parameter WEIGHT_0_5499 = 16'd-3403;
parameter WEIGHT_0_5500 = 16'd-2760;
parameter WEIGHT_0_5501 = 16'd1957;
parameter WEIGHT_0_5502 = 16'd2987;
parameter WEIGHT_0_5503 = 16'd7387;
parameter WEIGHT_0_5504 = 16'd-2530;
parameter WEIGHT_0_5505 = 16'd-683;
parameter WEIGHT_0_5506 = 16'd3875;
parameter WEIGHT_0_5507 = 16'd-8386;
parameter WEIGHT_0_5508 = 16'd-1537;
parameter WEIGHT_0_5509 = 16'd-2179;
parameter WEIGHT_0_5510 = 16'd-3139;
parameter WEIGHT_0_5511 = 16'd3382;
parameter WEIGHT_0_5512 = 16'd2247;
parameter WEIGHT_0_5513 = 16'd6463;
parameter WEIGHT_0_5514 = 16'd-8333;
parameter WEIGHT_0_5515 = 16'd996;
parameter WEIGHT_0_5516 = 16'd1538;
parameter WEIGHT_0_5517 = 16'd-8226;
parameter WEIGHT_0_5518 = 16'd977;
parameter WEIGHT_0_5519 = 16'd-2372;
parameter WEIGHT_0_5520 = 16'd-2312;
parameter WEIGHT_0_5521 = 16'd-81;
parameter WEIGHT_0_5522 = 16'd3332;
parameter WEIGHT_0_5523 = 16'd1523;
parameter WEIGHT_0_5524 = 16'd-4551;
parameter WEIGHT_0_5525 = 16'd3213;
parameter WEIGHT_0_5526 = 16'd1603;
parameter WEIGHT_0_5527 = 16'd-8228;
parameter WEIGHT_0_5528 = 16'd574;
parameter WEIGHT_0_5529 = 16'd-788;
parameter WEIGHT_0_5530 = 16'd362;
parameter WEIGHT_0_5531 = 16'd2663;
parameter WEIGHT_0_5532 = 16'd3945;
parameter WEIGHT_0_5533 = 16'd6199;
parameter WEIGHT_0_5534 = 16'd-4470;
parameter WEIGHT_0_5535 = 16'd1592;
parameter WEIGHT_0_5536 = 16'd-662;
parameter WEIGHT_0_5537 = 16'd-11355;
parameter WEIGHT_0_5538 = 16'd-320;
parameter WEIGHT_0_5539 = 16'd-6690;
parameter WEIGHT_0_5540 = 16'd12;
parameter WEIGHT_0_5541 = 16'd-3158;
parameter WEIGHT_0_5542 = 16'd5417;
parameter WEIGHT_0_5543 = 16'd1928;
parameter WEIGHT_0_5544 = 16'd-12330;
parameter WEIGHT_0_5545 = 16'd3220;
parameter WEIGHT_0_5546 = 16'd-2280;
parameter WEIGHT_0_5547 = 16'd-15848;
parameter WEIGHT_0_5548 = 16'd131;
parameter WEIGHT_0_5549 = 16'd-8751;
parameter WEIGHT_0_5550 = 16'd478;
parameter WEIGHT_0_5551 = 16'd-5258;
parameter WEIGHT_0_5552 = 16'd4258;
parameter WEIGHT_0_5553 = 16'd-653;
parameter WEIGHT_0_5554 = 16'd-11776;
parameter WEIGHT_0_5555 = 16'd3649;
parameter WEIGHT_0_5556 = 16'd-1513;
parameter WEIGHT_0_5557 = 16'd-16160;
parameter WEIGHT_0_5558 = 16'd462;
parameter WEIGHT_0_5559 = 16'd-12316;
parameter WEIGHT_0_5560 = 16'd-3585;
parameter WEIGHT_0_5561 = 16'd-1295;
parameter WEIGHT_0_5562 = 16'd7934;
parameter WEIGHT_0_5563 = 16'd-7282;
parameter WEIGHT_0_5564 = 16'd-12940;
parameter WEIGHT_0_5565 = 16'd5611;
parameter WEIGHT_0_5566 = 16'd-6127;
parameter WEIGHT_0_5567 = 16'd-6564;
parameter WEIGHT_0_5568 = 16'd-4301;
parameter WEIGHT_0_5569 = 16'd-7318;
parameter WEIGHT_0_5570 = 16'd-8413;
parameter WEIGHT_0_5571 = 16'd-1159;
parameter WEIGHT_0_5572 = 16'd14848;
parameter WEIGHT_0_5573 = 16'd-15337;
parameter WEIGHT_0_5574 = 16'd-12077;
parameter WEIGHT_0_5575 = 16'd-2847;
parameter WEIGHT_0_5576 = 16'd-6086;
parameter WEIGHT_0_5577 = 16'd-8229;
parameter WEIGHT_0_5578 = 16'd-18388;
parameter WEIGHT_0_5579 = 16'd-7624;
parameter WEIGHT_0_5580 = 16'd-7936;
parameter WEIGHT_0_5581 = 16'd1107;
parameter WEIGHT_0_5582 = 16'd9669;
parameter WEIGHT_0_5583 = 16'd-8660;
parameter WEIGHT_0_5584 = 16'd-2941;
parameter WEIGHT_0_5585 = 16'd-7939;
parameter WEIGHT_0_5586 = 16'd-9262;
parameter WEIGHT_0_5587 = 16'd-3534;
parameter WEIGHT_0_5588 = 16'd-7695;
parameter WEIGHT_0_5589 = 16'd-2556;
parameter WEIGHT_0_5590 = 16'd-5247;
parameter WEIGHT_0_5591 = 16'd4158;
parameter WEIGHT_0_5592 = 16'd4992;
parameter WEIGHT_0_5593 = 16'd-5231;
parameter WEIGHT_0_5594 = 16'd735;
parameter WEIGHT_0_5595 = 16'd-4955;
parameter WEIGHT_0_5596 = 16'd-1546;
parameter WEIGHT_0_5597 = 16'd1217;
parameter WEIGHT_0_5598 = 16'd-3487;
parameter WEIGHT_0_5599 = 16'd-1208;
parameter WEIGHT_0_5600 = 16'd-1491;
parameter WEIGHT_0_5601 = 16'd-1799;
parameter WEIGHT_0_5602 = 16'd-2085;
parameter WEIGHT_0_5603 = 16'd-2255;
parameter WEIGHT_0_5604 = 16'd-2343;
parameter WEIGHT_0_5605 = 16'd2463;
parameter WEIGHT_0_5606 = 16'd2833;
parameter WEIGHT_0_5607 = 16'd-110;
parameter WEIGHT_0_5608 = 16'd-2600;
parameter WEIGHT_0_5609 = 16'd2019;
parameter WEIGHT_0_5610 = 16'd-945;
parameter WEIGHT_0_5611 = 16'd-2339;
parameter WEIGHT_0_5612 = 16'd-5201;
parameter WEIGHT_0_5613 = 16'd-399;
parameter WEIGHT_0_5614 = 16'd-4607;
parameter WEIGHT_0_5615 = 16'd-8360;
parameter WEIGHT_0_5616 = 16'd-2094;
parameter WEIGHT_0_5617 = 16'd-363;
parameter WEIGHT_0_5618 = 16'd-4471;
parameter WEIGHT_0_5619 = 16'd-4413;
parameter WEIGHT_0_5620 = 16'd-3063;
parameter WEIGHT_0_5621 = 16'd-1701;
parameter WEIGHT_0_5622 = 16'd1569;
parameter WEIGHT_0_5623 = 16'd-1510;
parameter WEIGHT_0_5624 = 16'd-71;
parameter WEIGHT_0_5625 = 16'd-2049;
parameter WEIGHT_0_5626 = 16'd-4266;
parameter WEIGHT_0_5627 = 16'd-2704;
parameter WEIGHT_0_5628 = 16'd-9957;
parameter WEIGHT_0_5629 = 16'd-9189;
parameter WEIGHT_0_5630 = 16'd-7414;
parameter WEIGHT_0_5631 = 16'd-3618;
parameter WEIGHT_0_5632 = 16'd-2882;
parameter WEIGHT_0_5633 = 16'd10696;
parameter WEIGHT_0_5634 = 16'd-4877;
parameter WEIGHT_0_5635 = 16'd-1387;
parameter WEIGHT_0_5636 = 16'd-8774;
parameter WEIGHT_0_5637 = 16'd-9570;
parameter WEIGHT_0_5638 = 16'd-14314;
parameter WEIGHT_0_5639 = 16'd-12752;
parameter WEIGHT_0_5640 = 16'd-538;
parameter WEIGHT_0_5641 = 16'd-4962;
parameter WEIGHT_0_5642 = 16'd6030;
parameter WEIGHT_0_5643 = 16'd7175;
parameter WEIGHT_0_5644 = 16'd-7418;
parameter WEIGHT_0_5645 = 16'd-18;
parameter WEIGHT_0_5646 = 16'd-9221;
parameter WEIGHT_0_5647 = 16'd-14544;
parameter WEIGHT_0_5648 = 16'd-7943;
parameter WEIGHT_0_5649 = 16'd-7008;
parameter WEIGHT_0_5650 = 16'd3537;
parameter WEIGHT_0_5651 = 16'd-13254;
parameter WEIGHT_0_5652 = 16'd3850;
parameter WEIGHT_0_5653 = 16'd7212;
parameter WEIGHT_0_5654 = 16'd-8677;
parameter WEIGHT_0_5655 = 16'd2519;
parameter WEIGHT_0_5656 = 16'd-11163;
parameter WEIGHT_0_5657 = 16'd-10617;
parameter WEIGHT_0_5658 = 16'd-2573;
parameter WEIGHT_0_5659 = 16'd-4073;
parameter WEIGHT_0_5660 = 16'd2662;
parameter WEIGHT_0_5661 = 16'd-2921;
parameter WEIGHT_0_5662 = 16'd4231;
parameter WEIGHT_0_5663 = 16'd7132;
parameter WEIGHT_0_5664 = 16'd-12488;
parameter WEIGHT_0_5665 = 16'd5917;
parameter WEIGHT_0_5666 = 16'd-10053;
parameter WEIGHT_0_5667 = 16'd-12699;
parameter WEIGHT_0_5668 = 16'd-59;
parameter WEIGHT_0_5669 = 16'd-5201;
parameter WEIGHT_0_5670 = 16'd1444;
parameter WEIGHT_0_5671 = 16'd-2710;
parameter WEIGHT_0_5672 = 16'd6647;
parameter WEIGHT_0_5673 = 16'd1853;
parameter WEIGHT_0_5674 = 16'd-11993;
parameter WEIGHT_0_5675 = 16'd383;
parameter WEIGHT_0_5676 = 16'd-4315;
parameter WEIGHT_0_5677 = 16'd-15734;
parameter WEIGHT_0_5678 = 16'd4263;
parameter WEIGHT_0_5679 = 16'd-9395;
parameter WEIGHT_0_5680 = 16'd2430;
parameter WEIGHT_0_5681 = 16'd-972;
parameter WEIGHT_0_5682 = 16'd4448;
parameter WEIGHT_0_5683 = 16'd2819;
parameter WEIGHT_0_5684 = 16'd-15465;
parameter WEIGHT_0_5685 = 16'd5155;
parameter WEIGHT_0_5686 = 16'd-2288;
parameter WEIGHT_0_5687 = 16'd-11269;
parameter WEIGHT_0_5688 = 16'd1649;
parameter WEIGHT_0_5689 = 16'd-11126;
parameter WEIGHT_0_5690 = 16'd2537;
parameter WEIGHT_0_5691 = 16'd-5;
parameter WEIGHT_0_5692 = 16'd5337;
parameter WEIGHT_0_5693 = 16'd2164;
parameter WEIGHT_0_5694 = 16'd-12583;
parameter WEIGHT_0_5695 = 16'd4691;
parameter WEIGHT_0_5696 = 16'd1294;
parameter WEIGHT_0_5697 = 16'd-9107;
parameter WEIGHT_0_5698 = 16'd-1962;
parameter WEIGHT_0_5699 = 16'd-12898;
parameter WEIGHT_0_5700 = 16'd6375;
parameter WEIGHT_0_5701 = 16'd2011;
parameter WEIGHT_0_5702 = 16'd5092;
parameter WEIGHT_0_5703 = 16'd-4180;
parameter WEIGHT_0_5704 = 16'd-15759;
parameter WEIGHT_0_5705 = 16'd3095;
parameter WEIGHT_0_5706 = 16'd5872;
parameter WEIGHT_0_5707 = 16'd-9001;
parameter WEIGHT_0_5708 = 16'd-1218;
parameter WEIGHT_0_5709 = 16'd-14560;
parameter WEIGHT_0_5710 = 16'd6923;
parameter WEIGHT_0_5711 = 16'd2705;
parameter WEIGHT_0_5712 = 16'd5242;
parameter WEIGHT_0_5713 = 16'd-6667;
parameter WEIGHT_0_5714 = 16'd-7982;
parameter WEIGHT_0_5715 = 16'd5325;
parameter WEIGHT_0_5716 = 16'd7334;
parameter WEIGHT_0_5717 = 16'd-2661;
parameter WEIGHT_0_5718 = 16'd-4830;
parameter WEIGHT_0_5719 = 16'd-10935;
parameter WEIGHT_0_5720 = 16'd7600;
parameter WEIGHT_0_5721 = 16'd-730;
parameter WEIGHT_0_5722 = 16'd486;
parameter WEIGHT_0_5723 = 16'd-7558;
parameter WEIGHT_0_5724 = 16'd-8660;
parameter WEIGHT_0_5725 = 16'd-663;
parameter WEIGHT_0_5726 = 16'd9027;
parameter WEIGHT_0_5727 = 16'd-1539;
parameter WEIGHT_0_5728 = 16'd-4151;
parameter WEIGHT_0_5729 = 16'd-9753;
parameter WEIGHT_0_5730 = 16'd612;
parameter WEIGHT_0_5731 = 16'd-2622;
parameter WEIGHT_0_5732 = 16'd1391;
parameter WEIGHT_0_5733 = 16'd-4810;
parameter WEIGHT_0_5734 = 16'd-7565;
parameter WEIGHT_0_5735 = 16'd1882;
parameter WEIGHT_0_5736 = 16'd11610;
parameter WEIGHT_0_5737 = 16'd-621;
parameter WEIGHT_0_5738 = 16'd-3375;
parameter WEIGHT_0_5739 = 16'd-3672;
parameter WEIGHT_0_5740 = 16'd1674;
parameter WEIGHT_0_5741 = 16'd340;
parameter WEIGHT_0_5742 = 16'd1516;
parameter WEIGHT_0_5743 = 16'd1438;
parameter WEIGHT_0_5744 = 16'd144;
parameter WEIGHT_0_5745 = 16'd-565;
parameter WEIGHT_0_5746 = 16'd10502;
parameter WEIGHT_0_5747 = 16'd2657;
parameter WEIGHT_0_5748 = 16'd-3456;
parameter WEIGHT_0_5749 = 16'd-4524;
parameter WEIGHT_0_5750 = 16'd-2475;
parameter WEIGHT_0_5751 = 16'd-993;
parameter WEIGHT_0_5752 = 16'd1457;
parameter WEIGHT_0_5753 = 16'd2463;
parameter WEIGHT_0_5754 = 16'd-115;
parameter WEIGHT_0_5755 = 16'd376;
parameter WEIGHT_0_5756 = 16'd6561;
parameter WEIGHT_0_5757 = 16'd-2588;
parameter WEIGHT_0_5758 = 16'd346;
parameter WEIGHT_0_5759 = 16'd-5979;
parameter WEIGHT_0_5760 = 16'd1118;
parameter WEIGHT_0_5761 = 16'd4976;
parameter WEIGHT_0_5762 = 16'd1753;
parameter WEIGHT_0_5763 = 16'd4569;
parameter WEIGHT_0_5764 = 16'd1334;
parameter WEIGHT_0_5765 = 16'd408;
parameter WEIGHT_0_5766 = 16'd6999;
parameter WEIGHT_0_5767 = 16'd-5746;
parameter WEIGHT_0_5768 = 16'd-6257;
parameter WEIGHT_0_5769 = 16'd-3800;
parameter WEIGHT_0_5770 = 16'd-2286;
parameter WEIGHT_0_5771 = 16'd2604;
parameter WEIGHT_0_5772 = 16'd1682;
parameter WEIGHT_0_5773 = 16'd4141;
parameter WEIGHT_0_5774 = 16'd-1319;
parameter WEIGHT_0_5775 = 16'd3601;
parameter WEIGHT_0_5776 = 16'd3949;
parameter WEIGHT_0_5777 = 16'd-8177;
parameter WEIGHT_0_5778 = 16'd-482;
parameter WEIGHT_0_5779 = 16'd-5523;
parameter WEIGHT_0_5780 = 16'd-2081;
parameter WEIGHT_0_5781 = 16'd5973;
parameter WEIGHT_0_5782 = 16'd1120;
parameter WEIGHT_0_5783 = 16'd5387;
parameter WEIGHT_0_5784 = 16'd-3350;
parameter WEIGHT_0_5785 = 16'd4439;
parameter WEIGHT_0_5786 = 16'd2902;
parameter WEIGHT_0_5787 = 16'd-11295;
parameter WEIGHT_0_5788 = 16'd707;
parameter WEIGHT_0_5789 = 16'd-6681;
parameter WEIGHT_0_5790 = 16'd-2663;
parameter WEIGHT_0_5791 = 16'd5923;
parameter WEIGHT_0_5792 = 16'd2036;
parameter WEIGHT_0_5793 = 16'd4479;
parameter WEIGHT_0_5794 = 16'd-6465;
parameter WEIGHT_0_5795 = 16'd405;
parameter WEIGHT_0_5796 = 16'd2556;
parameter WEIGHT_0_5797 = 16'd-10934;
parameter WEIGHT_0_5798 = 16'd-839;
parameter WEIGHT_0_5799 = 16'd-1221;
parameter WEIGHT_0_5800 = 16'd-1314;
parameter WEIGHT_0_5801 = 16'd1328;
parameter WEIGHT_0_5802 = 16'd6068;
parameter WEIGHT_0_5803 = 16'd6241;
parameter WEIGHT_0_5804 = 16'd-4158;
parameter WEIGHT_0_5805 = 16'd143;
parameter WEIGHT_0_5806 = 16'd2514;
parameter WEIGHT_0_5807 = 16'd-16254;
parameter WEIGHT_0_5808 = 16'd214;
parameter WEIGHT_0_5809 = 16'd-3728;
parameter WEIGHT_0_5810 = 16'd709;
parameter WEIGHT_0_5811 = 16'd-773;
parameter WEIGHT_0_5812 = 16'd5395;
parameter WEIGHT_0_5813 = 16'd-47;
parameter WEIGHT_0_5814 = 16'd-3706;
parameter WEIGHT_0_5815 = 16'd1774;
parameter WEIGHT_0_5816 = 16'd-993;
parameter WEIGHT_0_5817 = 16'd-13542;
parameter WEIGHT_0_5818 = 16'd1916;
parameter WEIGHT_0_5819 = 16'd-9204;
parameter WEIGHT_0_5820 = 16'd-1882;
parameter WEIGHT_0_5821 = 16'd-183;
parameter WEIGHT_0_5822 = 16'd5635;
parameter WEIGHT_0_5823 = 16'd-2953;
parameter WEIGHT_0_5824 = 16'd-6976;
parameter WEIGHT_0_5825 = 16'd2799;
parameter WEIGHT_0_5826 = 16'd-3884;
parameter WEIGHT_0_5827 = 16'd-16994;
parameter WEIGHT_0_5828 = 16'd4453;
parameter WEIGHT_0_5829 = 16'd-8300;
parameter WEIGHT_0_5830 = 16'd-2180;
parameter WEIGHT_0_5831 = 16'd-6035;
parameter WEIGHT_0_5832 = 16'd4502;
parameter WEIGHT_0_5833 = 16'd-4489;
parameter WEIGHT_0_5834 = 16'd-11881;
parameter WEIGHT_0_5835 = 16'd2083;
parameter WEIGHT_0_5836 = 16'd-6851;
parameter WEIGHT_0_5837 = 16'd-14735;
parameter WEIGHT_0_5838 = 16'd4065;
parameter WEIGHT_0_5839 = 16'd-2450;
parameter WEIGHT_0_5840 = 16'd-7495;
parameter WEIGHT_0_5841 = 16'd451;
parameter WEIGHT_0_5842 = 16'd8327;
parameter WEIGHT_0_5843 = 16'd-5744;
parameter WEIGHT_0_5844 = 16'd-9555;
parameter WEIGHT_0_5845 = 16'd-1543;
parameter WEIGHT_0_5846 = 16'd-7111;
parameter WEIGHT_0_5847 = 16'd-5725;
parameter WEIGHT_0_5848 = 16'd-8413;
parameter WEIGHT_0_5849 = 16'd344;
parameter WEIGHT_0_5850 = 16'd-7746;
parameter WEIGHT_0_5851 = 16'd-436;
parameter WEIGHT_0_5852 = 16'd7592;
parameter WEIGHT_0_5853 = 16'd-16399;
parameter WEIGHT_0_5854 = 16'd-8118;
parameter WEIGHT_0_5855 = 16'd-1384;
parameter WEIGHT_0_5856 = 16'd-4171;
parameter WEIGHT_0_5857 = 16'd-9509;
parameter WEIGHT_0_5858 = 16'd-13871;
parameter WEIGHT_0_5859 = 16'd-168;
parameter WEIGHT_0_5860 = 16'd-1240;
parameter WEIGHT_0_5861 = 16'd726;
parameter WEIGHT_0_5862 = 16'd6652;
parameter WEIGHT_0_5863 = 16'd-4383;
parameter WEIGHT_0_5864 = 16'd-3272;
parameter WEIGHT_0_5865 = 16'd-3342;
parameter WEIGHT_0_5866 = 16'd-6105;
parameter WEIGHT_0_5867 = 16'd-3187;
parameter WEIGHT_0_5868 = 16'd-7172;
parameter WEIGHT_0_5869 = 16'd-1978;
parameter WEIGHT_0_5870 = 16'd-3011;
parameter WEIGHT_0_5871 = 16'd4163;
parameter WEIGHT_0_5872 = 16'd-5124;
parameter WEIGHT_0_5873 = 16'd-3402;
parameter WEIGHT_0_5874 = 16'd-3759;
parameter WEIGHT_0_5875 = 16'd3235;
parameter WEIGHT_0_5876 = 16'd-2640;
parameter WEIGHT_0_5877 = 16'd-2923;
parameter WEIGHT_0_5878 = 16'd-3063;
parameter WEIGHT_0_5879 = 16'd406;
parameter WEIGHT_0_5880 = 16'd-2138;
parameter WEIGHT_0_5881 = 16'd-348;
parameter WEIGHT_0_5882 = 16'd-46;
parameter WEIGHT_0_5883 = 16'd-2466;
parameter WEIGHT_0_5884 = 16'd994;
parameter WEIGHT_0_5885 = 16'd-1968;
parameter WEIGHT_0_5886 = 16'd-859;
parameter WEIGHT_0_5887 = 16'd-1696;
parameter WEIGHT_0_5888 = 16'd-3493;
parameter WEIGHT_0_5889 = 16'd-2203;
parameter WEIGHT_0_5890 = 16'd-4407;
parameter WEIGHT_0_5891 = 16'd2527;
parameter WEIGHT_0_5892 = 16'd1559;
parameter WEIGHT_0_5893 = 16'd1070;
parameter WEIGHT_0_5894 = 16'd-724;
parameter WEIGHT_0_5895 = 16'd-8579;
parameter WEIGHT_0_5896 = 16'd-420;
parameter WEIGHT_0_5897 = 16'd-3856;
parameter WEIGHT_0_5898 = 16'd-2847;
parameter WEIGHT_0_5899 = 16'd-1302;
parameter WEIGHT_0_5900 = 16'd-3739;
parameter WEIGHT_0_5901 = 16'd-2856;
parameter WEIGHT_0_5902 = 16'd-693;
parameter WEIGHT_0_5903 = 16'd4527;
parameter WEIGHT_0_5904 = 16'd-1439;
parameter WEIGHT_0_5905 = 16'd-4987;
parameter WEIGHT_0_5906 = 16'd-3303;
parameter WEIGHT_0_5907 = 16'd-7393;
parameter WEIGHT_0_5908 = 16'd-10502;
parameter WEIGHT_0_5909 = 16'd-7852;
parameter WEIGHT_0_5910 = 16'd-5575;
parameter WEIGHT_0_5911 = 16'd-3039;
parameter WEIGHT_0_5912 = 16'd3100;
parameter WEIGHT_0_5913 = 16'd10320;
parameter WEIGHT_0_5914 = 16'd-6077;
parameter WEIGHT_0_5915 = 16'd-376;
parameter WEIGHT_0_5916 = 16'd-9779;
parameter WEIGHT_0_5917 = 16'd-14370;
parameter WEIGHT_0_5918 = 16'd-14051;
parameter WEIGHT_0_5919 = 16'd-13639;
parameter WEIGHT_0_5920 = 16'd-5772;
parameter WEIGHT_0_5921 = 16'd2757;
parameter WEIGHT_0_5922 = 16'd602;
parameter WEIGHT_0_5923 = 16'd6403;
parameter WEIGHT_0_5924 = 16'd-8908;
parameter WEIGHT_0_5925 = 16'd2853;
parameter WEIGHT_0_5926 = 16'd-14505;
parameter WEIGHT_0_5927 = 16'd-8668;
parameter WEIGHT_0_5928 = 16'd-8406;
parameter WEIGHT_0_5929 = 16'd-5062;
parameter WEIGHT_0_5930 = 16'd1024;
parameter WEIGHT_0_5931 = 16'd2795;
parameter WEIGHT_0_5932 = 16'd870;
parameter WEIGHT_0_5933 = 16'd3704;
parameter WEIGHT_0_5934 = 16'd-7769;
parameter WEIGHT_0_5935 = 16'd1106;
parameter WEIGHT_0_5936 = 16'd-15467;
parameter WEIGHT_0_5937 = 16'd-10271;
parameter WEIGHT_0_5938 = 16'd-348;
parameter WEIGHT_0_5939 = 16'd-2520;
parameter WEIGHT_0_5940 = 16'd-1750;
parameter WEIGHT_0_5941 = 16'd5315;
parameter WEIGHT_0_5942 = 16'd657;
parameter WEIGHT_0_5943 = 16'd3753;
parameter WEIGHT_0_5944 = 16'd-15274;
parameter WEIGHT_0_5945 = 16'd-423;
parameter WEIGHT_0_5946 = 16'd-12354;
parameter WEIGHT_0_5947 = 16'd-8535;
parameter WEIGHT_0_5948 = 16'd1624;
parameter WEIGHT_0_5949 = 16'd-7277;
parameter WEIGHT_0_5950 = 16'd558;
parameter WEIGHT_0_5951 = 16'd469;
parameter WEIGHT_0_5952 = 16'd4204;
parameter WEIGHT_0_5953 = 16'd3236;
parameter WEIGHT_0_5954 = 16'd-15652;
parameter WEIGHT_0_5955 = 16'd666;
parameter WEIGHT_0_5956 = 16'd-6482;
parameter WEIGHT_0_5957 = 16'd-7332;
parameter WEIGHT_0_5958 = 16'd3597;
parameter WEIGHT_0_5959 = 16'd-6237;
parameter WEIGHT_0_5960 = 16'd602;
parameter WEIGHT_0_5961 = 16'd2071;
parameter WEIGHT_0_5962 = 16'd337;
parameter WEIGHT_0_5963 = 16'd578;
parameter WEIGHT_0_5964 = 16'd-9559;
parameter WEIGHT_0_5965 = 16'd5186;
parameter WEIGHT_0_5966 = 16'd-2775;
parameter WEIGHT_0_5967 = 16'd-5061;
parameter WEIGHT_0_5968 = 16'd507;
parameter WEIGHT_0_5969 = 16'd-4113;
parameter WEIGHT_0_5970 = 16'd2185;
parameter WEIGHT_0_5971 = 16'd86;
parameter WEIGHT_0_5972 = 16'd2715;
parameter WEIGHT_0_5973 = 16'd-1903;
parameter WEIGHT_0_5974 = 16'd-10383;
parameter WEIGHT_0_5975 = 16'd1538;
parameter WEIGHT_0_5976 = 16'd-1007;
parameter WEIGHT_0_5977 = 16'd-5025;
parameter WEIGHT_0_5978 = 16'd-619;
parameter WEIGHT_0_5979 = 16'd-8130;
parameter WEIGHT_0_5980 = 16'd3668;
parameter WEIGHT_0_5981 = 16'd-64;
parameter WEIGHT_0_5982 = 16'd2154;
parameter WEIGHT_0_5983 = 16'd-705;
parameter WEIGHT_0_5984 = 16'd-7758;
parameter WEIGHT_0_5985 = 16'd2921;
parameter WEIGHT_0_5986 = 16'd2862;
parameter WEIGHT_0_5987 = 16'd-5612;
parameter WEIGHT_0_5988 = 16'd-3028;
parameter WEIGHT_0_5989 = 16'd-6828;
parameter WEIGHT_0_5990 = 16'd5427;
parameter WEIGHT_0_5991 = 16'd-3147;
parameter WEIGHT_0_5992 = 16'd4622;
parameter WEIGHT_0_5993 = 16'd-4039;
parameter WEIGHT_0_5994 = 16'd-3797;
parameter WEIGHT_0_5995 = 16'd1339;
parameter WEIGHT_0_5996 = 16'd6072;
parameter WEIGHT_0_5997 = 16'd-2200;
parameter WEIGHT_0_5998 = 16'd-567;
parameter WEIGHT_0_5999 = 16'd-9919;
parameter WEIGHT_0_6000 = 16'd7181;
parameter WEIGHT_0_6001 = 16'd-7358;
parameter WEIGHT_0_6002 = 16'd1288;
parameter WEIGHT_0_6003 = 16'd-3022;
parameter WEIGHT_0_6004 = 16'd-7059;
parameter WEIGHT_0_6005 = 16'd1193;
parameter WEIGHT_0_6006 = 16'd11427;
parameter WEIGHT_0_6007 = 16'd500;
parameter WEIGHT_0_6008 = 16'd-2042;
parameter WEIGHT_0_6009 = 16'd-7412;
parameter WEIGHT_0_6010 = 16'd345;
parameter WEIGHT_0_6011 = 16'd-3753;
parameter WEIGHT_0_6012 = 16'd914;
parameter WEIGHT_0_6013 = 16'd-1797;
parameter WEIGHT_0_6014 = 16'd-8662;
parameter WEIGHT_0_6015 = 16'd14;
parameter WEIGHT_0_6016 = 16'd9816;
parameter WEIGHT_0_6017 = 16'd588;
parameter WEIGHT_0_6018 = 16'd2756;
parameter WEIGHT_0_6019 = 16'd-5717;
parameter WEIGHT_0_6020 = 16'd-222;
parameter WEIGHT_0_6021 = 16'd-1875;
parameter WEIGHT_0_6022 = 16'd-2916;
parameter WEIGHT_0_6023 = 16'd-1130;
parameter WEIGHT_0_6024 = 16'd-2277;
parameter WEIGHT_0_6025 = 16'd2740;
parameter WEIGHT_0_6026 = 16'd11491;
parameter WEIGHT_0_6027 = 16'd-1245;
parameter WEIGHT_0_6028 = 16'd214;
parameter WEIGHT_0_6029 = 16'd-4768;
parameter WEIGHT_0_6030 = 16'd-56;
parameter WEIGHT_0_6031 = 16'd282;
parameter WEIGHT_0_6032 = 16'd-1414;
parameter WEIGHT_0_6033 = 16'd1559;
parameter WEIGHT_0_6034 = 16'd-2547;
parameter WEIGHT_0_6035 = 16'd2817;
parameter WEIGHT_0_6036 = 16'd8951;
parameter WEIGHT_0_6037 = 16'd-2197;
parameter WEIGHT_0_6038 = 16'd704;
parameter WEIGHT_0_6039 = 16'd-4348;
parameter WEIGHT_0_6040 = 16'd-1224;
parameter WEIGHT_0_6041 = 16'd2631;
parameter WEIGHT_0_6042 = 16'd1853;
parameter WEIGHT_0_6043 = 16'd2479;
parameter WEIGHT_0_6044 = 16'd-1843;
parameter WEIGHT_0_6045 = 16'd1875;
parameter WEIGHT_0_6046 = 16'd5476;
parameter WEIGHT_0_6047 = 16'd-2387;
parameter WEIGHT_0_6048 = 16'd-1487;
parameter WEIGHT_0_6049 = 16'd-1746;
parameter WEIGHT_0_6050 = 16'd-3172;
parameter WEIGHT_0_6051 = 16'd5396;
parameter WEIGHT_0_6052 = 16'd2155;
parameter WEIGHT_0_6053 = 16'd1540;
parameter WEIGHT_0_6054 = 16'd-1027;
parameter WEIGHT_0_6055 = 16'd3510;
parameter WEIGHT_0_6056 = 16'd5992;
parameter WEIGHT_0_6057 = 16'd-9459;
parameter WEIGHT_0_6058 = 16'd-3095;
parameter WEIGHT_0_6059 = 16'd-6753;
parameter WEIGHT_0_6060 = 16'd-5108;
parameter WEIGHT_0_6061 = 16'd5284;
parameter WEIGHT_0_6062 = 16'd6686;
parameter WEIGHT_0_6063 = 16'd4283;
parameter WEIGHT_0_6064 = 16'd-4497;
parameter WEIGHT_0_6065 = 16'd-486;
parameter WEIGHT_0_6066 = 16'd4771;
parameter WEIGHT_0_6067 = 16'd-10477;
parameter WEIGHT_0_6068 = 16'd-765;
parameter WEIGHT_0_6069 = 16'd-6596;
parameter WEIGHT_0_6070 = 16'd-6603;
parameter WEIGHT_0_6071 = 16'd525;
parameter WEIGHT_0_6072 = 16'd6662;
parameter WEIGHT_0_6073 = 16'd3320;
parameter WEIGHT_0_6074 = 16'd-2534;
parameter WEIGHT_0_6075 = 16'd-13;
parameter WEIGHT_0_6076 = 16'd409;
parameter WEIGHT_0_6077 = 16'd-10449;
parameter WEIGHT_0_6078 = 16'd-696;
parameter WEIGHT_0_6079 = 16'd-7407;
parameter WEIGHT_0_6080 = 16'd-3088;
parameter WEIGHT_0_6081 = 16'd4639;
parameter WEIGHT_0_6082 = 16'd2718;
parameter WEIGHT_0_6083 = 16'd2549;
parameter WEIGHT_0_6084 = 16'd-2779;
parameter WEIGHT_0_6085 = 16'd1709;
parameter WEIGHT_0_6086 = 16'd315;
parameter WEIGHT_0_6087 = 16'd-12371;
parameter WEIGHT_0_6088 = 16'd2746;
parameter WEIGHT_0_6089 = 16'd-1776;
parameter WEIGHT_0_6090 = 16'd-2221;
parameter WEIGHT_0_6091 = 16'd-1232;
parameter WEIGHT_0_6092 = 16'd2139;
parameter WEIGHT_0_6093 = 16'd-3106;
parameter WEIGHT_0_6094 = 16'd-2784;
parameter WEIGHT_0_6095 = 16'd6083;
parameter WEIGHT_0_6096 = 16'd-3619;
parameter WEIGHT_0_6097 = 16'd-14445;
parameter WEIGHT_0_6098 = 16'd-1150;
parameter WEIGHT_0_6099 = 16'd-6433;
parameter WEIGHT_0_6100 = 16'd-269;
parameter WEIGHT_0_6101 = 16'd-5124;
parameter WEIGHT_0_6102 = 16'd6615;
parameter WEIGHT_0_6103 = 16'd-4844;
parameter WEIGHT_0_6104 = 16'd-4169;
parameter WEIGHT_0_6105 = 16'd7654;
parameter WEIGHT_0_6106 = 16'd-5604;
parameter WEIGHT_0_6107 = 16'd-16955;
parameter WEIGHT_0_6108 = 16'd3608;
parameter WEIGHT_0_6109 = 16'd-1834;
parameter WEIGHT_0_6110 = 16'd-2987;
parameter WEIGHT_0_6111 = 16'd-8522;
parameter WEIGHT_0_6112 = 16'd8290;
parameter WEIGHT_0_6113 = 16'd-7527;
parameter WEIGHT_0_6114 = 16'd-2537;
parameter WEIGHT_0_6115 = 16'd6345;
parameter WEIGHT_0_6116 = 16'd-5214;
parameter WEIGHT_0_6117 = 16'd-16115;
parameter WEIGHT_0_6118 = 16'd-2837;
parameter WEIGHT_0_6119 = 16'd-3294;
parameter WEIGHT_0_6120 = 16'd-5859;
parameter WEIGHT_0_6121 = 16'd1347;
parameter WEIGHT_0_6122 = 16'd10461;
parameter WEIGHT_0_6123 = 16'd-13185;
parameter WEIGHT_0_6124 = 16'd-7596;
parameter WEIGHT_0_6125 = 16'd266;
parameter WEIGHT_0_6126 = 16'd-7861;
parameter WEIGHT_0_6127 = 16'd-6369;
parameter WEIGHT_0_6128 = 16'd-8933;
parameter WEIGHT_0_6129 = 16'd4268;
parameter WEIGHT_0_6130 = 16'd-8255;
parameter WEIGHT_0_6131 = 16'd-448;
parameter WEIGHT_0_6132 = 16'd8060;
parameter WEIGHT_0_6133 = 16'd-9599;
parameter WEIGHT_0_6134 = 16'd-9536;
parameter WEIGHT_0_6135 = 16'd562;
parameter WEIGHT_0_6136 = 16'd-3561;
parameter WEIGHT_0_6137 = 16'd-1630;
parameter WEIGHT_0_6138 = 16'd-9126;
parameter WEIGHT_0_6139 = 16'd1177;
parameter WEIGHT_0_6140 = 16'd587;
parameter WEIGHT_0_6141 = 16'd-1978;
parameter WEIGHT_0_6142 = 16'd1014;
parameter WEIGHT_0_6143 = 16'd-5840;
parameter WEIGHT_0_6144 = 16'd-3121;
parameter WEIGHT_0_6145 = 16'd1955;
parameter WEIGHT_0_6146 = 16'd-2672;
parameter WEIGHT_0_6147 = 16'd-2453;
parameter WEIGHT_0_6148 = 16'd-8352;
parameter WEIGHT_0_6149 = 16'd-6663;
parameter WEIGHT_0_6150 = 16'd-1104;
parameter WEIGHT_0_6151 = 16'd-2130;
parameter WEIGHT_0_6152 = 16'd-3100;
parameter WEIGHT_0_6153 = 16'd-2757;
parameter WEIGHT_0_6154 = 16'd-2392;
parameter WEIGHT_0_6155 = 16'd-461;
parameter WEIGHT_0_6156 = 16'd-2146;
parameter WEIGHT_0_6157 = 16'd699;
parameter WEIGHT_0_6158 = 16'd-3344;
parameter WEIGHT_0_6159 = 16'd-847;
parameter WEIGHT_0_6160 = 16'd-687;
parameter WEIGHT_0_6161 = 16'd4586;
parameter WEIGHT_0_6162 = 16'd-2374;
parameter WEIGHT_0_6163 = 16'd-4037;
parameter WEIGHT_0_6164 = 16'd1512;
parameter WEIGHT_0_6165 = 16'd1792;
parameter WEIGHT_0_6166 = 16'd282;
parameter WEIGHT_0_6167 = 16'd1334;
parameter WEIGHT_0_6168 = 16'd-4501;
parameter WEIGHT_0_6169 = 16'd-7;
parameter WEIGHT_0_6170 = 16'd651;
parameter WEIGHT_0_6171 = 16'd-370;
parameter WEIGHT_0_6172 = 16'd-1104;
parameter WEIGHT_0_6173 = 16'd-711;
parameter WEIGHT_0_6174 = 16'd-1176;
parameter WEIGHT_0_6175 = 16'd-2363;
parameter WEIGHT_0_6176 = 16'd-2900;
parameter WEIGHT_0_6177 = 16'd-1789;
parameter WEIGHT_0_6178 = 16'd-1701;
parameter WEIGHT_0_6179 = 16'd-1733;
parameter WEIGHT_0_6180 = 16'd-5315;
parameter WEIGHT_0_6181 = 16'd-1475;
parameter WEIGHT_0_6182 = 16'd-1365;
parameter WEIGHT_0_6183 = 16'd4172;
parameter WEIGHT_0_6184 = 16'd-156;
parameter WEIGHT_0_6185 = 16'd-9758;
parameter WEIGHT_0_6186 = 16'd-2523;
parameter WEIGHT_0_6187 = 16'd-8020;
parameter WEIGHT_0_6188 = 16'd-6747;
parameter WEIGHT_0_6189 = 16'd-7052;
parameter WEIGHT_0_6190 = 16'd-7441;
parameter WEIGHT_0_6191 = 16'd-2968;
parameter WEIGHT_0_6192 = 16'd2853;
parameter WEIGHT_0_6193 = 16'd9118;
parameter WEIGHT_0_6194 = 16'd-6628;
parameter WEIGHT_0_6195 = 16'd-336;
parameter WEIGHT_0_6196 = 16'd-4110;
parameter WEIGHT_0_6197 = 16'd-10595;
parameter WEIGHT_0_6198 = 16'd-7069;
parameter WEIGHT_0_6199 = 16'd-2890;
parameter WEIGHT_0_6200 = 16'd-9864;
parameter WEIGHT_0_6201 = 16'd2256;
parameter WEIGHT_0_6202 = 16'd2490;
parameter WEIGHT_0_6203 = 16'd4052;
parameter WEIGHT_0_6204 = 16'd-8987;
parameter WEIGHT_0_6205 = 16'd1488;
parameter WEIGHT_0_6206 = 16'd-16043;
parameter WEIGHT_0_6207 = 16'd-3653;
parameter WEIGHT_0_6208 = 16'd-7449;
parameter WEIGHT_0_6209 = 16'd-6233;
parameter WEIGHT_0_6210 = 16'd906;
parameter WEIGHT_0_6211 = 16'd14889;
parameter WEIGHT_0_6212 = 16'd2294;
parameter WEIGHT_0_6213 = 16'd4560;
parameter WEIGHT_0_6214 = 16'd-15940;
parameter WEIGHT_0_6215 = 16'd-182;
parameter WEIGHT_0_6216 = 16'd-16462;
parameter WEIGHT_0_6217 = 16'd-1622;
parameter WEIGHT_0_6218 = 16'd-4719;
parameter WEIGHT_0_6219 = 16'd-9353;
parameter WEIGHT_0_6220 = 16'd-299;
parameter WEIGHT_0_6221 = 16'd9571;
parameter WEIGHT_0_6222 = 16'd6166;
parameter WEIGHT_0_6223 = 16'd2678;
parameter WEIGHT_0_6224 = 16'd-9678;
parameter WEIGHT_0_6225 = 16'd-2344;
parameter WEIGHT_0_6226 = 16'd-20102;
parameter WEIGHT_0_6227 = 16'd-4165;
parameter WEIGHT_0_6228 = 16'd656;
parameter WEIGHT_0_6229 = 16'd-7451;
parameter WEIGHT_0_6230 = 16'd1868;
parameter WEIGHT_0_6231 = 16'd5844;
parameter WEIGHT_0_6232 = 16'd2806;
parameter WEIGHT_0_6233 = 16'd2255;
parameter WEIGHT_0_6234 = 16'd-9890;
parameter WEIGHT_0_6235 = 16'd-2446;
parameter WEIGHT_0_6236 = 16'd-12221;
parameter WEIGHT_0_6237 = 16'd2650;
parameter WEIGHT_0_6238 = 16'd556;
parameter WEIGHT_0_6239 = 16'd-8299;
parameter WEIGHT_0_6240 = 16'd1201;
parameter WEIGHT_0_6241 = 16'd-589;
parameter WEIGHT_0_6242 = 16'd6166;
parameter WEIGHT_0_6243 = 16'd-1197;
parameter WEIGHT_0_6244 = 16'd-6300;
parameter WEIGHT_0_6245 = 16'd48;
parameter WEIGHT_0_6246 = 16'd-3330;
parameter WEIGHT_0_6247 = 16'd-1769;
parameter WEIGHT_0_6248 = 16'd-334;
parameter WEIGHT_0_6249 = 16'd-1449;
parameter WEIGHT_0_6250 = 16'd3164;
parameter WEIGHT_0_6251 = 16'd3214;
parameter WEIGHT_0_6252 = 16'd5738;
parameter WEIGHT_0_6253 = 16'd734;
parameter WEIGHT_0_6254 = 16'd-8167;
parameter WEIGHT_0_6255 = 16'd-776;
parameter WEIGHT_0_6256 = 16'd-4128;
parameter WEIGHT_0_6257 = 16'd-3485;
parameter WEIGHT_0_6258 = 16'd-2495;
parameter WEIGHT_0_6259 = 16'd-1433;
parameter WEIGHT_0_6260 = 16'd2076;
parameter WEIGHT_0_6261 = 16'd-943;
parameter WEIGHT_0_6262 = 16'd4104;
parameter WEIGHT_0_6263 = 16'd1496;
parameter WEIGHT_0_6264 = 16'd-2258;
parameter WEIGHT_0_6265 = 16'd1779;
parameter WEIGHT_0_6266 = 16'd1301;
parameter WEIGHT_0_6267 = 16'd-3868;
parameter WEIGHT_0_6268 = 16'd-1169;
parameter WEIGHT_0_6269 = 16'd631;
parameter WEIGHT_0_6270 = 16'd7075;
parameter WEIGHT_0_6271 = 16'd-6000;
parameter WEIGHT_0_6272 = 16'd4036;
parameter WEIGHT_0_6273 = 16'd-110;
parameter WEIGHT_0_6274 = 16'd-6213;
parameter WEIGHT_0_6275 = 16'd2840;
parameter WEIGHT_0_6276 = 16'd-819;
parameter WEIGHT_0_6277 = 16'd-3537;
parameter WEIGHT_0_6278 = 16'd1793;
parameter WEIGHT_0_6279 = 16'd-2196;
parameter WEIGHT_0_6280 = 16'd3911;
parameter WEIGHT_0_6281 = 16'd-8361;
parameter WEIGHT_0_6282 = 16'd-18;
parameter WEIGHT_0_6283 = 16'd-337;
parameter WEIGHT_0_6284 = 16'd-3056;
parameter WEIGHT_0_6285 = 16'd5435;
parameter WEIGHT_0_6286 = 16'd4086;
parameter WEIGHT_0_6287 = 16'd-903;
parameter WEIGHT_0_6288 = 16'd4482;
parameter WEIGHT_0_6289 = 16'd-3329;
parameter WEIGHT_0_6290 = 16'd8178;
parameter WEIGHT_0_6291 = 16'd-12436;
parameter WEIGHT_0_6292 = 16'd-2018;
parameter WEIGHT_0_6293 = 16'd-2563;
parameter WEIGHT_0_6294 = 16'd-7125;
parameter WEIGHT_0_6295 = 16'd3474;
parameter WEIGHT_0_6296 = 16'd4094;
parameter WEIGHT_0_6297 = 16'd-5818;
parameter WEIGHT_0_6298 = 16'd4650;
parameter WEIGHT_0_6299 = 16'd-2726;
parameter WEIGHT_0_6300 = 16'd5179;
parameter WEIGHT_0_6301 = 16'd-1231;
parameter WEIGHT_0_6302 = 16'd-2093;
parameter WEIGHT_0_6303 = 16'd-1898;
parameter WEIGHT_0_6304 = 16'd-3740;
parameter WEIGHT_0_6305 = 16'd2328;
parameter WEIGHT_0_6306 = 16'd-115;
parameter WEIGHT_0_6307 = 16'd468;
parameter WEIGHT_0_6308 = 16'd2451;
parameter WEIGHT_0_6309 = 16'd-1786;
parameter WEIGHT_0_6310 = 16'd2968;
parameter WEIGHT_0_6311 = 16'd433;
parameter WEIGHT_0_6312 = 16'd-2701;
parameter WEIGHT_0_6313 = 16'd1501;
parameter WEIGHT_0_6314 = 16'd-1175;
parameter WEIGHT_0_6315 = 16'd2079;
parameter WEIGHT_0_6316 = 16'd846;
parameter WEIGHT_0_6317 = 16'd-1896;
parameter WEIGHT_0_6318 = 16'd1350;
parameter WEIGHT_0_6319 = 16'd-6316;
parameter WEIGHT_0_6320 = 16'd1659;
parameter WEIGHT_0_6321 = 16'd1646;
parameter WEIGHT_0_6322 = 16'd-2231;
parameter WEIGHT_0_6323 = 16'd4393;
parameter WEIGHT_0_6324 = 16'd-1419;
parameter WEIGHT_0_6325 = 16'd4274;
parameter WEIGHT_0_6326 = 16'd2479;
parameter WEIGHT_0_6327 = 16'd-4013;
parameter WEIGHT_0_6328 = 16'd1620;
parameter WEIGHT_0_6329 = 16'd-3512;
parameter WEIGHT_0_6330 = 16'd-3085;
parameter WEIGHT_0_6331 = 16'd5932;
parameter WEIGHT_0_6332 = 16'd207;
parameter WEIGHT_0_6333 = 16'd1249;
parameter WEIGHT_0_6334 = 16'd19;
parameter WEIGHT_0_6335 = 16'd-816;
parameter WEIGHT_0_6336 = 16'd-2611;
parameter WEIGHT_0_6337 = 16'd-4687;
parameter WEIGHT_0_6338 = 16'd-1657;
parameter WEIGHT_0_6339 = 16'd-7448;
parameter WEIGHT_0_6340 = 16'd-4147;
parameter WEIGHT_0_6341 = 16'd4982;
parameter WEIGHT_0_6342 = 16'd6410;
parameter WEIGHT_0_6343 = 16'd2015;
parameter WEIGHT_0_6344 = 16'd1189;
parameter WEIGHT_0_6345 = 16'd3474;
parameter WEIGHT_0_6346 = 16'd-2954;
parameter WEIGHT_0_6347 = 16'd-9762;
parameter WEIGHT_0_6348 = 16'd1636;
parameter WEIGHT_0_6349 = 16'd-5755;
parameter WEIGHT_0_6350 = 16'd-1545;
parameter WEIGHT_0_6351 = 16'd4566;
parameter WEIGHT_0_6352 = 16'd6637;
parameter WEIGHT_0_6353 = 16'd2252;
parameter WEIGHT_0_6354 = 16'd4392;
parameter WEIGHT_0_6355 = 16'd1825;
parameter WEIGHT_0_6356 = 16'd-508;
parameter WEIGHT_0_6357 = 16'd-8427;
parameter WEIGHT_0_6358 = 16'd-2141;
parameter WEIGHT_0_6359 = 16'd-5369;
parameter WEIGHT_0_6360 = 16'd-2021;
parameter WEIGHT_0_6361 = 16'd4396;
parameter WEIGHT_0_6362 = 16'd4663;
parameter WEIGHT_0_6363 = 16'd2013;
parameter WEIGHT_0_6364 = 16'd2124;
parameter WEIGHT_0_6365 = 16'd5279;
parameter WEIGHT_0_6366 = 16'd-4876;
parameter WEIGHT_0_6367 = 16'd-13761;
parameter WEIGHT_0_6368 = 16'd-509;
parameter WEIGHT_0_6369 = 16'd-4800;
parameter WEIGHT_0_6370 = 16'd-5614;
parameter WEIGHT_0_6371 = 16'd-1780;
parameter WEIGHT_0_6372 = 16'd5482;
parameter WEIGHT_0_6373 = 16'd-1689;
parameter WEIGHT_0_6374 = 16'd3291;
parameter WEIGHT_0_6375 = 16'd1635;
parameter WEIGHT_0_6376 = 16'd-4365;
parameter WEIGHT_0_6377 = 16'd-13882;
parameter WEIGHT_0_6378 = 16'd1682;
parameter WEIGHT_0_6379 = 16'd-1500;
parameter WEIGHT_0_6380 = 16'd-3832;
parameter WEIGHT_0_6381 = 16'd-7460;
parameter WEIGHT_0_6382 = 16'd6359;
parameter WEIGHT_0_6383 = 16'd-3370;
parameter WEIGHT_0_6384 = 16'd-2526;
parameter WEIGHT_0_6385 = 16'd3001;
parameter WEIGHT_0_6386 = 16'd-9076;
parameter WEIGHT_0_6387 = 16'd-14265;
parameter WEIGHT_0_6388 = 16'd-582;
parameter WEIGHT_0_6389 = 16'd1615;
parameter WEIGHT_0_6390 = 16'd-1609;
parameter WEIGHT_0_6391 = 16'd-3620;
parameter WEIGHT_0_6392 = 16'd2601;
parameter WEIGHT_0_6393 = 16'd-7525;
parameter WEIGHT_0_6394 = 16'd-2557;
parameter WEIGHT_0_6395 = 16'd4338;
parameter WEIGHT_0_6396 = 16'd-8842;
parameter WEIGHT_0_6397 = 16'd-14258;
parameter WEIGHT_0_6398 = 16'd-1975;
parameter WEIGHT_0_6399 = 16'd1445;
parameter WEIGHT_0_6400 = 16'd-6946;
parameter WEIGHT_0_6401 = 16'd-2432;
parameter WEIGHT_0_6402 = 16'd8879;
parameter WEIGHT_0_6403 = 16'd-11507;
parameter WEIGHT_0_6404 = 16'd-254;
parameter WEIGHT_0_6405 = 16'd3308;
parameter WEIGHT_0_6406 = 16'd-9148;
parameter WEIGHT_0_6407 = 16'd-6754;
parameter WEIGHT_0_6408 = 16'd-6518;
parameter WEIGHT_0_6409 = 16'd4815;
parameter WEIGHT_0_6410 = 16'd-1423;
parameter WEIGHT_0_6411 = 16'd-1081;
parameter WEIGHT_0_6412 = 16'd5948;
parameter WEIGHT_0_6413 = 16'd-7969;
parameter WEIGHT_0_6414 = 16'd-4781;
parameter WEIGHT_0_6415 = 16'd2104;
parameter WEIGHT_0_6416 = 16'd-8557;
parameter WEIGHT_0_6417 = 16'd-4767;
parameter WEIGHT_0_6418 = 16'd-9743;
parameter WEIGHT_0_6419 = 16'd1714;
parameter WEIGHT_0_6420 = 16'd1911;
parameter WEIGHT_0_6421 = 16'd2874;
parameter WEIGHT_0_6422 = 16'd-2329;
parameter WEIGHT_0_6423 = 16'd746;
parameter WEIGHT_0_6424 = 16'd3692;
parameter WEIGHT_0_6425 = 16'd19;
parameter WEIGHT_0_6426 = 16'd3069;
parameter WEIGHT_0_6427 = 16'd-6929;
parameter WEIGHT_0_6428 = 16'd-4963;
parameter WEIGHT_0_6429 = 16'd-8517;
parameter WEIGHT_0_6430 = 16'd-831;
parameter WEIGHT_0_6431 = 16'd1107;
parameter WEIGHT_0_6432 = 16'd1522;
parameter WEIGHT_0_6433 = 16'd791;
parameter WEIGHT_0_6434 = 16'd2429;
parameter WEIGHT_0_6435 = 16'd1941;
parameter WEIGHT_0_6436 = 16'd1342;
parameter WEIGHT_0_6437 = 16'd-3217;
parameter WEIGHT_0_6438 = 16'd-3290;
parameter WEIGHT_0_6439 = 16'd-2777;
parameter WEIGHT_0_6440 = 16'd-863;
parameter WEIGHT_0_6441 = 16'd753;
parameter WEIGHT_0_6442 = 16'd1002;
parameter WEIGHT_0_6443 = 16'd2533;
parameter WEIGHT_0_6444 = 16'd2759;
parameter WEIGHT_0_6445 = 16'd-650;
parameter WEIGHT_0_6446 = 16'd-2686;
parameter WEIGHT_0_6447 = 16'd-1012;
parameter WEIGHT_0_6448 = 16'd-646;
parameter WEIGHT_0_6449 = 16'd1636;
parameter WEIGHT_0_6450 = 16'd-1791;
parameter WEIGHT_0_6451 = 16'd-556;
parameter WEIGHT_0_6452 = 16'd-1457;
parameter WEIGHT_0_6453 = 16'd-2688;
parameter WEIGHT_0_6454 = 16'd996;
parameter WEIGHT_0_6455 = 16'd1302;
parameter WEIGHT_0_6456 = 16'd-1920;
parameter WEIGHT_0_6457 = 16'd-724;
parameter WEIGHT_0_6458 = 16'd2634;
parameter WEIGHT_0_6459 = 16'd-1730;
parameter WEIGHT_0_6460 = 16'd-1097;
parameter WEIGHT_0_6461 = 16'd-3633;
parameter WEIGHT_0_6462 = 16'd-2361;
parameter WEIGHT_0_6463 = 16'd7969;
parameter WEIGHT_0_6464 = 16'd-1314;
parameter WEIGHT_0_6465 = 16'd-2950;
parameter WEIGHT_0_6466 = 16'd-3100;
parameter WEIGHT_0_6467 = 16'd-3226;
parameter WEIGHT_0_6468 = 16'd-5190;
parameter WEIGHT_0_6469 = 16'd-7629;
parameter WEIGHT_0_6470 = 16'd-7222;
parameter WEIGHT_0_6471 = 16'd-6193;
parameter WEIGHT_0_6472 = 16'd-2336;
parameter WEIGHT_0_6473 = 16'd10818;
parameter WEIGHT_0_6474 = 16'd-4420;
parameter WEIGHT_0_6475 = 16'd2917;
parameter WEIGHT_0_6476 = 16'd-5345;
parameter WEIGHT_0_6477 = 16'd-10536;
parameter WEIGHT_0_6478 = 16'd-8674;
parameter WEIGHT_0_6479 = 16'd-3728;
parameter WEIGHT_0_6480 = 16'd-12966;
parameter WEIGHT_0_6481 = 16'd-2156;
parameter WEIGHT_0_6482 = 16'd-3108;
parameter WEIGHT_0_6483 = 16'd7706;
parameter WEIGHT_0_6484 = 16'd-11777;
parameter WEIGHT_0_6485 = 16'd3839;
parameter WEIGHT_0_6486 = 16'd-7731;
parameter WEIGHT_0_6487 = 16'd2367;
parameter WEIGHT_0_6488 = 16'd-12133;
parameter WEIGHT_0_6489 = 16'd-5935;
parameter WEIGHT_0_6490 = 16'd-6843;
parameter WEIGHT_0_6491 = 16'd6325;
parameter WEIGHT_0_6492 = 16'd-548;
parameter WEIGHT_0_6493 = 16'd9356;
parameter WEIGHT_0_6494 = 16'd-10880;
parameter WEIGHT_0_6495 = 16'd2320;
parameter WEIGHT_0_6496 = 16'd-11025;
parameter WEIGHT_0_6497 = 16'd5241;
parameter WEIGHT_0_6498 = 16'd-10991;
parameter WEIGHT_0_6499 = 16'd-5612;
parameter WEIGHT_0_6500 = 16'd230;
parameter WEIGHT_0_6501 = 16'd5958;
parameter WEIGHT_0_6502 = 16'd-783;
parameter WEIGHT_0_6503 = 16'd6827;
parameter WEIGHT_0_6504 = 16'd-7067;
parameter WEIGHT_0_6505 = 16'd-3648;
parameter WEIGHT_0_6506 = 16'd-15713;
parameter WEIGHT_0_6507 = 16'd5080;
parameter WEIGHT_0_6508 = 16'd-9743;
parameter WEIGHT_0_6509 = 16'd-3243;
parameter WEIGHT_0_6510 = 16'd1811;
parameter WEIGHT_0_6511 = 16'd3022;
parameter WEIGHT_0_6512 = 16'd119;
parameter WEIGHT_0_6513 = 16'd3299;
parameter WEIGHT_0_6514 = 16'd-1961;
parameter WEIGHT_0_6515 = 16'd-3521;
parameter WEIGHT_0_6516 = 16'd-17812;
parameter WEIGHT_0_6517 = 16'd4906;
parameter WEIGHT_0_6518 = 16'd-3216;
parameter WEIGHT_0_6519 = 16'd-5675;
parameter WEIGHT_0_6520 = 16'd1394;
parameter WEIGHT_0_6521 = 16'd-1162;
parameter WEIGHT_0_6522 = 16'd167;
parameter WEIGHT_0_6523 = 16'd3411;
parameter WEIGHT_0_6524 = 16'd-3177;
parameter WEIGHT_0_6525 = 16'd-501;
parameter WEIGHT_0_6526 = 16'd-13302;
parameter WEIGHT_0_6527 = 16'd-3176;
parameter WEIGHT_0_6528 = 16'd-1535;
parameter WEIGHT_0_6529 = 16'd2236;
parameter WEIGHT_0_6530 = 16'd3521;
parameter WEIGHT_0_6531 = 16'd-1777;
parameter WEIGHT_0_6532 = 16'd2695;
parameter WEIGHT_0_6533 = 16'd2979;
parameter WEIGHT_0_6534 = 16'd-2765;
parameter WEIGHT_0_6535 = 16'd1733;
parameter WEIGHT_0_6536 = 16'd-9210;
parameter WEIGHT_0_6537 = 16'd1027;
parameter WEIGHT_0_6538 = 16'd1701;
parameter WEIGHT_0_6539 = 16'd-2243;
parameter WEIGHT_0_6540 = 16'd7984;
parameter WEIGHT_0_6541 = 16'd-4338;
parameter WEIGHT_0_6542 = 16'd-2791;
parameter WEIGHT_0_6543 = 16'd4303;
parameter WEIGHT_0_6544 = 16'd-3636;
parameter WEIGHT_0_6545 = 16'd4632;
parameter WEIGHT_0_6546 = 16'd-10166;
parameter WEIGHT_0_6547 = 16'd-3346;
parameter WEIGHT_0_6548 = 16'd1198;
parameter WEIGHT_0_6549 = 16'd-2686;
parameter WEIGHT_0_6550 = 16'd6919;
parameter WEIGHT_0_6551 = 16'd-7978;
parameter WEIGHT_0_6552 = 16'd1600;
parameter WEIGHT_0_6553 = 16'd756;
parameter WEIGHT_0_6554 = 16'd-2100;
parameter WEIGHT_0_6555 = 16'd3183;
parameter WEIGHT_0_6556 = 16'd-9879;
parameter WEIGHT_0_6557 = 16'd-2924;
parameter WEIGHT_0_6558 = 16'd2135;
parameter WEIGHT_0_6559 = 16'd-1464;
parameter WEIGHT_0_6560 = 16'd5781;
parameter WEIGHT_0_6561 = 16'd-6302;
parameter WEIGHT_0_6562 = 16'd-2106;
parameter WEIGHT_0_6563 = 16'd1576;
parameter WEIGHT_0_6564 = 16'd-4853;
parameter WEIGHT_0_6565 = 16'd1407;
parameter WEIGHT_0_6566 = 16'd-6730;
parameter WEIGHT_0_6567 = 16'd-4625;
parameter WEIGHT_0_6568 = 16'd4095;
parameter WEIGHT_0_6569 = 16'd-4261;
parameter WEIGHT_0_6570 = 16'd7216;
parameter WEIGHT_0_6571 = 16'd-6468;
parameter WEIGHT_0_6572 = 16'd-2809;
parameter WEIGHT_0_6573 = 16'd1214;
parameter WEIGHT_0_6574 = 16'd-5914;
parameter WEIGHT_0_6575 = 16'd3145;
parameter WEIGHT_0_6576 = 16'd-6995;
parameter WEIGHT_0_6577 = 16'd-1239;
parameter WEIGHT_0_6578 = 16'd7500;
parameter WEIGHT_0_6579 = 16'd-6370;
parameter WEIGHT_0_6580 = 16'd5536;
parameter WEIGHT_0_6581 = 16'd-3945;
parameter WEIGHT_0_6582 = 16'd-4359;
parameter WEIGHT_0_6583 = 16'd549;
parameter WEIGHT_0_6584 = 16'd-3888;
parameter WEIGHT_0_6585 = 16'd2529;
parameter WEIGHT_0_6586 = 16'd-2752;
parameter WEIGHT_0_6587 = 16'd-1243;
parameter WEIGHT_0_6588 = 16'd8208;
parameter WEIGHT_0_6589 = 16'd-3007;
parameter WEIGHT_0_6590 = 16'd1842;
parameter WEIGHT_0_6591 = 16'd1555;
parameter WEIGHT_0_6592 = 16'd-744;
parameter WEIGHT_0_6593 = 16'd-941;
parameter WEIGHT_0_6594 = 16'd-3496;
parameter WEIGHT_0_6595 = 16'd2328;
parameter WEIGHT_0_6596 = 16'd-2470;
parameter WEIGHT_0_6597 = 16'd2127;
parameter WEIGHT_0_6598 = 16'd5893;
parameter WEIGHT_0_6599 = 16'd-6780;
parameter WEIGHT_0_6600 = 16'd1367;
parameter WEIGHT_0_6601 = 16'd2521;
parameter WEIGHT_0_6602 = 16'd-3009;
parameter WEIGHT_0_6603 = 16'd-1576;
parameter WEIGHT_0_6604 = 16'd1840;
parameter WEIGHT_0_6605 = 16'd2811;
parameter WEIGHT_0_6606 = 16'd-4114;
parameter WEIGHT_0_6607 = 16'd1946;
parameter WEIGHT_0_6608 = 16'd5594;
parameter WEIGHT_0_6609 = 16'd-3093;
parameter WEIGHT_0_6610 = 16'd-1895;
parameter WEIGHT_0_6611 = 16'd10666;
parameter WEIGHT_0_6612 = 16'd-289;
parameter WEIGHT_0_6613 = 16'd3935;
parameter WEIGHT_0_6614 = 16'd3766;
parameter WEIGHT_0_6615 = 16'd359;
parameter WEIGHT_0_6616 = 16'd-5383;
parameter WEIGHT_0_6617 = 16'd-1539;
parameter WEIGHT_0_6618 = 16'd1146;
parameter WEIGHT_0_6619 = 16'd-2102;
parameter WEIGHT_0_6620 = 16'd-6108;
parameter WEIGHT_0_6621 = 16'd1318;
parameter WEIGHT_0_6622 = 16'd3753;
parameter WEIGHT_0_6623 = 16'd1465;
parameter WEIGHT_0_6624 = 16'd2818;
parameter WEIGHT_0_6625 = 16'd-1668;
parameter WEIGHT_0_6626 = 16'd-5302;
parameter WEIGHT_0_6627 = 16'd-5346;
parameter WEIGHT_0_6628 = 16'd3979;
parameter WEIGHT_0_6629 = 16'd-3199;
parameter WEIGHT_0_6630 = 16'd-6674;
parameter WEIGHT_0_6631 = 16'd1104;
parameter WEIGHT_0_6632 = 16'd4927;
parameter WEIGHT_0_6633 = 16'd960;
parameter WEIGHT_0_6634 = 16'd5926;
parameter WEIGHT_0_6635 = 16'd-646;
parameter WEIGHT_0_6636 = 16'd-2068;
parameter WEIGHT_0_6637 = 16'd-9065;
parameter WEIGHT_0_6638 = 16'd-605;
parameter WEIGHT_0_6639 = 16'd692;
parameter WEIGHT_0_6640 = 16'd-10432;
parameter WEIGHT_0_6641 = 16'd-3863;
parameter WEIGHT_0_6642 = 16'd7195;
parameter WEIGHT_0_6643 = 16'd-4855;
parameter WEIGHT_0_6644 = 16'd2789;
parameter WEIGHT_0_6645 = 16'd-478;
parameter WEIGHT_0_6646 = 16'd-4791;
parameter WEIGHT_0_6647 = 16'd-11721;
parameter WEIGHT_0_6648 = 16'd1679;
parameter WEIGHT_0_6649 = 16'd-931;
parameter WEIGHT_0_6650 = 16'd-6013;
parameter WEIGHT_0_6651 = 16'd-3933;
parameter WEIGHT_0_6652 = 16'd3166;
parameter WEIGHT_0_6653 = 16'd-7753;
parameter WEIGHT_0_6654 = 16'd6245;
parameter WEIGHT_0_6655 = 16'd1068;
parameter WEIGHT_0_6656 = 16'd-8734;
parameter WEIGHT_0_6657 = 16'd-13865;
parameter WEIGHT_0_6658 = 16'd-19;
parameter WEIGHT_0_6659 = 16'd3600;
parameter WEIGHT_0_6660 = 16'd-5277;
parameter WEIGHT_0_6661 = 16'd-5182;
parameter WEIGHT_0_6662 = 16'd6791;
parameter WEIGHT_0_6663 = 16'd-5932;
parameter WEIGHT_0_6664 = 16'd633;
parameter WEIGHT_0_6665 = 16'd2093;
parameter WEIGHT_0_6666 = 16'd-9163;
parameter WEIGHT_0_6667 = 16'd-10757;
parameter WEIGHT_0_6668 = 16'd1458;
parameter WEIGHT_0_6669 = 16'd6184;
parameter WEIGHT_0_6670 = 16'd-5839;
parameter WEIGHT_0_6671 = 16'd-10055;
parameter WEIGHT_0_6672 = 16'd5894;
parameter WEIGHT_0_6673 = 16'd-9089;
parameter WEIGHT_0_6674 = 16'd-5320;
parameter WEIGHT_0_6675 = 16'd3592;
parameter WEIGHT_0_6676 = 16'd-12629;
parameter WEIGHT_0_6677 = 16'd-17405;
parameter WEIGHT_0_6678 = 16'd3292;
parameter WEIGHT_0_6679 = 16'd8096;
parameter WEIGHT_0_6680 = 16'd-2949;
parameter WEIGHT_0_6681 = 16'd-6309;
parameter WEIGHT_0_6682 = 16'd5967;
parameter WEIGHT_0_6683 = 16'd-5335;
parameter WEIGHT_0_6684 = 16'd-6106;
parameter WEIGHT_0_6685 = 16'd3341;
parameter WEIGHT_0_6686 = 16'd-9581;
parameter WEIGHT_0_6687 = 16'd-3875;
parameter WEIGHT_0_6688 = 16'd-3322;
parameter WEIGHT_0_6689 = 16'd4769;
parameter WEIGHT_0_6690 = 16'd-2549;
parameter WEIGHT_0_6691 = 16'd19;
parameter WEIGHT_0_6692 = 16'd4927;
parameter WEIGHT_0_6693 = 16'd-5508;
parameter WEIGHT_0_6694 = 16'd-3530;
parameter WEIGHT_0_6695 = 16'd-656;
parameter WEIGHT_0_6696 = 16'd-4788;
parameter WEIGHT_0_6697 = 16'd-5438;
parameter WEIGHT_0_6698 = 16'd-6824;
parameter WEIGHT_0_6699 = 16'd-2010;
parameter WEIGHT_0_6700 = 16'd-5682;
parameter WEIGHT_0_6701 = 16'd2929;
parameter WEIGHT_0_6702 = 16'd-5311;
parameter WEIGHT_0_6703 = 16'd1718;
parameter WEIGHT_0_6704 = 16'd2181;
parameter WEIGHT_0_6705 = 16'd3059;
parameter WEIGHT_0_6706 = 16'd-83;
parameter WEIGHT_0_6707 = 16'd-5876;
parameter WEIGHT_0_6708 = 16'd-5049;
parameter WEIGHT_0_6709 = 16'd-4066;
parameter WEIGHT_0_6710 = 16'd-1;
parameter WEIGHT_0_6711 = 16'd-874;
parameter WEIGHT_0_6712 = 16'd2190;
parameter WEIGHT_0_6713 = 16'd-1357;
parameter WEIGHT_0_6714 = 16'd519;
parameter WEIGHT_0_6715 = 16'd1720;
parameter WEIGHT_0_6716 = 16'd-1981;
parameter WEIGHT_0_6717 = 16'd572;
parameter WEIGHT_0_6718 = 16'd-1845;
parameter WEIGHT_0_6719 = 16'd-1079;
parameter WEIGHT_0_6720 = 16'd-2120;
parameter WEIGHT_0_6721 = 16'd2019;
parameter WEIGHT_0_6722 = 16'd2800;
parameter WEIGHT_0_6723 = 16'd-179;
parameter WEIGHT_0_6724 = 16'd1112;
parameter WEIGHT_0_6725 = 16'd111;
parameter WEIGHT_0_6726 = 16'd251;
parameter WEIGHT_0_6727 = 16'd-2744;
parameter WEIGHT_0_6728 = 16'd2225;
parameter WEIGHT_0_6729 = 16'd2544;
parameter WEIGHT_0_6730 = 16'd-2085;
parameter WEIGHT_0_6731 = 16'd2467;
parameter WEIGHT_0_6732 = 16'd1524;
parameter WEIGHT_0_6733 = 16'd2232;
parameter WEIGHT_0_6734 = 16'd1625;
parameter WEIGHT_0_6735 = 16'd-1292;
parameter WEIGHT_0_6736 = 16'd-2661;
parameter WEIGHT_0_6737 = 16'd-284;
parameter WEIGHT_0_6738 = 16'd-557;
parameter WEIGHT_0_6739 = 16'd344;
parameter WEIGHT_0_6740 = 16'd-2309;
parameter WEIGHT_0_6741 = 16'd-173;
parameter WEIGHT_0_6742 = 16'd-6568;
parameter WEIGHT_0_6743 = 16'd3947;
parameter WEIGHT_0_6744 = 16'd-2080;
parameter WEIGHT_0_6745 = 16'd-3891;
parameter WEIGHT_0_6746 = 16'd1034;
parameter WEIGHT_0_6747 = 16'd497;
parameter WEIGHT_0_6748 = 16'd-2661;
parameter WEIGHT_0_6749 = 16'd-4576;
parameter WEIGHT_0_6750 = 16'd-3914;
parameter WEIGHT_0_6751 = 16'd-5011;
parameter WEIGHT_0_6752 = 16'd-11015;
parameter WEIGHT_0_6753 = 16'd6059;
parameter WEIGHT_0_6754 = 16'd-4324;
parameter WEIGHT_0_6755 = 16'd-429;
parameter WEIGHT_0_6756 = 16'd-475;
parameter WEIGHT_0_6757 = 16'd-336;
parameter WEIGHT_0_6758 = 16'd-4107;
parameter WEIGHT_0_6759 = 16'd-8814;
parameter WEIGHT_0_6760 = 16'd-6727;
parameter WEIGHT_0_6761 = 16'd-6769;
parameter WEIGHT_0_6762 = 16'd-7991;
parameter WEIGHT_0_6763 = 16'd9259;
parameter WEIGHT_0_6764 = 16'd-8687;
parameter WEIGHT_0_6765 = 16'd-1112;
parameter WEIGHT_0_6766 = 16'd-3342;
parameter WEIGHT_0_6767 = 16'd5603;
parameter WEIGHT_0_6768 = 16'd-14571;
parameter WEIGHT_0_6769 = 16'd-2240;
parameter WEIGHT_0_6770 = 16'd-6664;
parameter WEIGHT_0_6771 = 16'd187;
parameter WEIGHT_0_6772 = 16'd-13112;
parameter WEIGHT_0_6773 = 16'd7581;
parameter WEIGHT_0_6774 = 16'd-6546;
parameter WEIGHT_0_6775 = 16'd-1086;
parameter WEIGHT_0_6776 = 16'd-10169;
parameter WEIGHT_0_6777 = 16'd11484;
parameter WEIGHT_0_6778 = 16'd-19423;
parameter WEIGHT_0_6779 = 16'd107;
parameter WEIGHT_0_6780 = 16'd-7020;
parameter WEIGHT_0_6781 = 16'd-289;
parameter WEIGHT_0_6782 = 16'd-13961;
parameter WEIGHT_0_6783 = 16'd9470;
parameter WEIGHT_0_6784 = 16'd-3297;
parameter WEIGHT_0_6785 = 16'd-289;
parameter WEIGHT_0_6786 = 16'd-13174;
parameter WEIGHT_0_6787 = 16'd11370;
parameter WEIGHT_0_6788 = 16'd-12627;
parameter WEIGHT_0_6789 = 16'd-496;
parameter WEIGHT_0_6790 = 16'd-8657;
parameter WEIGHT_0_6791 = 16'd-3161;
parameter WEIGHT_0_6792 = 16'd-8715;
parameter WEIGHT_0_6793 = 16'd11648;
parameter WEIGHT_0_6794 = 16'd-5313;
parameter WEIGHT_0_6795 = 16'd-2436;
parameter WEIGHT_0_6796 = 16'd-13279;
parameter WEIGHT_0_6797 = 16'd8380;
parameter WEIGHT_0_6798 = 16'd-7411;
parameter WEIGHT_0_6799 = 16'd5765;
parameter WEIGHT_0_6800 = 16'd-1800;
parameter WEIGHT_0_6801 = 16'd-5389;
parameter WEIGHT_0_6802 = 16'd-8685;
parameter WEIGHT_0_6803 = 16'd7765;
parameter WEIGHT_0_6804 = 16'd-2184;
parameter WEIGHT_0_6805 = 16'd522;
parameter WEIGHT_0_6806 = 16'd-14481;
parameter WEIGHT_0_6807 = 16'd8113;
parameter WEIGHT_0_6808 = 16'd-3256;
parameter WEIGHT_0_6809 = 16'd2254;
parameter WEIGHT_0_6810 = 16'd-5089;
parameter WEIGHT_0_6811 = 16'd-5472;
parameter WEIGHT_0_6812 = 16'd-7044;
parameter WEIGHT_0_6813 = 16'd4310;
parameter WEIGHT_0_6814 = 16'd-1893;
parameter WEIGHT_0_6815 = 16'd2949;
parameter WEIGHT_0_6816 = 16'd-17079;
parameter WEIGHT_0_6817 = 16'd1032;
parameter WEIGHT_0_6818 = 16'd-1034;
parameter WEIGHT_0_6819 = 16'd-623;
parameter WEIGHT_0_6820 = 16'd-965;
parameter WEIGHT_0_6821 = 16'd-8079;
parameter WEIGHT_0_6822 = 16'd-8826;
parameter WEIGHT_0_6823 = 16'd6520;
parameter WEIGHT_0_6824 = 16'd-2517;
parameter WEIGHT_0_6825 = 16'd4698;
parameter WEIGHT_0_6826 = 16'd-21875;
parameter WEIGHT_0_6827 = 16'd2907;
parameter WEIGHT_0_6828 = 16'd1393;
parameter WEIGHT_0_6829 = 16'd-118;
parameter WEIGHT_0_6830 = 16'd-3202;
parameter WEIGHT_0_6831 = 16'd-7684;
parameter WEIGHT_0_6832 = 16'd-6894;
parameter WEIGHT_0_6833 = 16'd7509;
parameter WEIGHT_0_6834 = 16'd-2143;
parameter WEIGHT_0_6835 = 16'd2456;
parameter WEIGHT_0_6836 = 16'd-19219;
parameter WEIGHT_0_6837 = 16'd2290;
parameter WEIGHT_0_6838 = 16'd390;
parameter WEIGHT_0_6839 = 16'd-1586;
parameter WEIGHT_0_6840 = 16'd4105;
parameter WEIGHT_0_6841 = 16'd-10164;
parameter WEIGHT_0_6842 = 16'd-1529;
parameter WEIGHT_0_6843 = 16'd4911;
parameter WEIGHT_0_6844 = 16'd-4505;
parameter WEIGHT_0_6845 = 16'd3724;
parameter WEIGHT_0_6846 = 16'd-13414;
parameter WEIGHT_0_6847 = 16'd2014;
parameter WEIGHT_0_6848 = 16'd2265;
parameter WEIGHT_0_6849 = 16'd-2649;
parameter WEIGHT_0_6850 = 16'd1621;
parameter WEIGHT_0_6851 = 16'd-8565;
parameter WEIGHT_0_6852 = 16'd-4033;
parameter WEIGHT_0_6853 = 16'd6299;
parameter WEIGHT_0_6854 = 16'd-3195;
parameter WEIGHT_0_6855 = 16'd8203;
parameter WEIGHT_0_6856 = 16'd-16725;
parameter WEIGHT_0_6857 = 16'd3724;
parameter WEIGHT_0_6858 = 16'd5976;
parameter WEIGHT_0_6859 = 16'd-3920;
parameter WEIGHT_0_6860 = 16'd-439;
parameter WEIGHT_0_6861 = 16'd-10644;
parameter WEIGHT_0_6862 = 16'd-444;
parameter WEIGHT_0_6863 = 16'd5312;
parameter WEIGHT_0_6864 = 16'd-3612;
parameter WEIGHT_0_6865 = 16'd3631;
parameter WEIGHT_0_6866 = 16'd-12092;
parameter WEIGHT_0_6867 = 16'd3758;
parameter WEIGHT_0_6868 = 16'd1991;
parameter WEIGHT_0_6869 = 16'd-5578;
parameter WEIGHT_0_6870 = 16'd1062;
parameter WEIGHT_0_6871 = 16'd-8097;
parameter WEIGHT_0_6872 = 16'd-2850;
parameter WEIGHT_0_6873 = 16'd2875;
parameter WEIGHT_0_6874 = 16'd-4929;
parameter WEIGHT_0_6875 = 16'd5712;
parameter WEIGHT_0_6876 = 16'd-12255;
parameter WEIGHT_0_6877 = 16'd2147;
parameter WEIGHT_0_6878 = 16'd4956;
parameter WEIGHT_0_6879 = 16'd-4017;
parameter WEIGHT_0_6880 = 16'd-5261;
parameter WEIGHT_0_6881 = 16'd-8239;
parameter WEIGHT_0_6882 = 16'd-3172;
parameter WEIGHT_0_6883 = 16'd1970;
parameter WEIGHT_0_6884 = 16'd-238;
parameter WEIGHT_0_6885 = 16'd2929;
parameter WEIGHT_0_6886 = 16'd-12729;
parameter WEIGHT_0_6887 = 16'd160;
parameter WEIGHT_0_6888 = 16'd6456;
parameter WEIGHT_0_6889 = 16'd53;
parameter WEIGHT_0_6890 = 16'd-3956;
parameter WEIGHT_0_6891 = 16'd-3304;
parameter WEIGHT_0_6892 = 16'd-169;
parameter WEIGHT_0_6893 = 16'd1336;
parameter WEIGHT_0_6894 = 16'd-2540;
parameter WEIGHT_0_6895 = 16'd1881;
parameter WEIGHT_0_6896 = 16'd-10774;
parameter WEIGHT_0_6897 = 16'd-1801;
parameter WEIGHT_0_6898 = 16'd1370;
parameter WEIGHT_0_6899 = 16'd2025;
parameter WEIGHT_0_6900 = 16'd-10964;
parameter WEIGHT_0_6901 = 16'd2534;
parameter WEIGHT_0_6902 = 16'd4059;
parameter WEIGHT_0_6903 = 16'd-2242;
parameter WEIGHT_0_6904 = 16'd957;
parameter WEIGHT_0_6905 = 16'd3983;
parameter WEIGHT_0_6906 = 16'd-10384;
parameter WEIGHT_0_6907 = 16'd-5729;
parameter WEIGHT_0_6908 = 16'd5182;
parameter WEIGHT_0_6909 = 16'd379;
parameter WEIGHT_0_6910 = 16'd-12456;
parameter WEIGHT_0_6911 = 16'd-1797;
parameter WEIGHT_0_6912 = 16'd-717;
parameter WEIGHT_0_6913 = 16'd-6827;
parameter WEIGHT_0_6914 = 16'd1273;
parameter WEIGHT_0_6915 = 16'd912;
parameter WEIGHT_0_6916 = 16'd-16536;
parameter WEIGHT_0_6917 = 16'd-5757;
parameter WEIGHT_0_6918 = 16'd5354;
parameter WEIGHT_0_6919 = 16'd5885;
parameter WEIGHT_0_6920 = 16'd-12245;
parameter WEIGHT_0_6921 = 16'd-1596;
parameter WEIGHT_0_6922 = 16'd-3524;
parameter WEIGHT_0_6923 = 16'd-5160;
parameter WEIGHT_0_6924 = 16'd-760;
parameter WEIGHT_0_6925 = 16'd1243;
parameter WEIGHT_0_6926 = 16'd-15874;
parameter WEIGHT_0_6927 = 16'd-5437;
parameter WEIGHT_0_6928 = 16'd2152;
parameter WEIGHT_0_6929 = 16'd5433;
parameter WEIGHT_0_6930 = 16'd-11666;
parameter WEIGHT_0_6931 = 16'd-3578;
parameter WEIGHT_0_6932 = 16'd2988;
parameter WEIGHT_0_6933 = 16'd-6442;
parameter WEIGHT_0_6934 = 16'd-886;
parameter WEIGHT_0_6935 = 16'd-542;
parameter WEIGHT_0_6936 = 16'd-16167;
parameter WEIGHT_0_6937 = 16'd-7572;
parameter WEIGHT_0_6938 = 16'd-4847;
parameter WEIGHT_0_6939 = 16'd9020;
parameter WEIGHT_0_6940 = 16'd-9222;
parameter WEIGHT_0_6941 = 16'd-4189;
parameter WEIGHT_0_6942 = 16'd791;
parameter WEIGHT_0_6943 = 16'd-7367;
parameter WEIGHT_0_6944 = 16'd-2602;
parameter WEIGHT_0_6945 = 16'd3925;
parameter WEIGHT_0_6946 = 16'd-9717;
parameter WEIGHT_0_6947 = 16'd-9339;
parameter WEIGHT_0_6948 = 16'd-5355;
parameter WEIGHT_0_6949 = 16'd10397;
parameter WEIGHT_0_6950 = 16'd-6710;
parameter WEIGHT_0_6951 = 16'd-8743;
parameter WEIGHT_0_6952 = 16'd174;
parameter WEIGHT_0_6953 = 16'd-6321;
parameter WEIGHT_0_6954 = 16'd-2034;
parameter WEIGHT_0_6955 = 16'd2538;
parameter WEIGHT_0_6956 = 16'd-8999;
parameter WEIGHT_0_6957 = 16'd-14851;
parameter WEIGHT_0_6958 = 16'd-3098;
parameter WEIGHT_0_6959 = 16'd5019;
parameter WEIGHT_0_6960 = 16'd-4493;
parameter WEIGHT_0_6961 = 16'd-3118;
parameter WEIGHT_0_6962 = 16'd7351;
parameter WEIGHT_0_6963 = 16'd-6020;
parameter WEIGHT_0_6964 = 16'd-5196;
parameter WEIGHT_0_6965 = 16'd1205;
parameter WEIGHT_0_6966 = 16'd-2215;
parameter WEIGHT_0_6967 = 16'd-9957;
parameter WEIGHT_0_6968 = 16'd-11414;
parameter WEIGHT_0_6969 = 16'd677;
parameter WEIGHT_0_6970 = 16'd-4822;
parameter WEIGHT_0_6971 = 16'd-289;
parameter WEIGHT_0_6972 = 16'd5537;
parameter WEIGHT_0_6973 = 16'd-3035;
parameter WEIGHT_0_6974 = 16'd-646;
parameter WEIGHT_0_6975 = 16'd-7138;
parameter WEIGHT_0_6976 = 16'd-5334;
parameter WEIGHT_0_6977 = 16'd-7627;
parameter WEIGHT_0_6978 = 16'd-9714;
parameter WEIGHT_0_6979 = 16'd-4128;
parameter WEIGHT_0_6980 = 16'd-3355;
parameter WEIGHT_0_6981 = 16'd4061;
parameter WEIGHT_0_6982 = 16'd1347;
parameter WEIGHT_0_6983 = 16'd-5363;
parameter WEIGHT_0_6984 = 16'd792;
parameter WEIGHT_0_6985 = 16'd-4971;
parameter WEIGHT_0_6986 = 16'd-4588;
parameter WEIGHT_0_6987 = 16'd-1307;
parameter WEIGHT_0_6988 = 16'd-4908;
parameter WEIGHT_0_6989 = 16'd-107;
parameter WEIGHT_0_6990 = 16'd-694;
parameter WEIGHT_0_6991 = 16'd2376;
parameter WEIGHT_0_6992 = 16'd-2066;
parameter WEIGHT_0_6993 = 16'd-2711;
parameter WEIGHT_0_6994 = 16'd-2518;
parameter WEIGHT_0_6995 = 16'd-594;
parameter WEIGHT_0_6996 = 16'd-1755;
parameter WEIGHT_0_6997 = 16'd2211;
parameter WEIGHT_0_6998 = 16'd-2346;
parameter WEIGHT_0_6999 = 16'd2800;
parameter WEIGHT_0_7000 = 16'd-2231;
parameter WEIGHT_0_7001 = 16'd535;
parameter WEIGHT_0_7002 = 16'd-1262;
parameter WEIGHT_0_7003 = 16'd953;
parameter WEIGHT_0_7004 = 16'd1887;
parameter WEIGHT_0_7005 = 16'd2246;
parameter WEIGHT_0_7006 = 16'd2115;
parameter WEIGHT_0_7007 = 16'd-969;
parameter WEIGHT_0_7008 = 16'd-459;
parameter WEIGHT_0_7009 = 16'd-1087;
parameter WEIGHT_0_7010 = 16'd1281;
parameter WEIGHT_0_7011 = 16'd1391;
parameter WEIGHT_0_7012 = 16'd-697;
parameter WEIGHT_0_7013 = 16'd-593;
parameter WEIGHT_0_7014 = 16'd-2534;
parameter WEIGHT_0_7015 = 16'd846;
parameter WEIGHT_0_7016 = 16'd809;
parameter WEIGHT_0_7017 = 16'd2332;
parameter WEIGHT_0_7018 = 16'd2127;
parameter WEIGHT_0_7019 = 16'd-389;
parameter WEIGHT_0_7020 = 16'd-4464;
parameter WEIGHT_0_7021 = 16'd126;
parameter WEIGHT_0_7022 = 16'd-1854;
parameter WEIGHT_0_7023 = 16'd3348;
parameter WEIGHT_0_7024 = 16'd-443;
parameter WEIGHT_0_7025 = 16'd1193;
parameter WEIGHT_0_7026 = 16'd1940;
parameter WEIGHT_0_7027 = 16'd-6509;
parameter WEIGHT_0_7028 = 16'd-3316;
parameter WEIGHT_0_7029 = 16'd1068;
parameter WEIGHT_0_7030 = 16'd-3226;
parameter WEIGHT_0_7031 = 16'd-2109;
parameter WEIGHT_0_7032 = 16'd-4661;
parameter WEIGHT_0_7033 = 16'd-2403;
parameter WEIGHT_0_7034 = 16'd1055;
parameter WEIGHT_0_7035 = 16'd2983;
parameter WEIGHT_0_7036 = 16'd-644;
parameter WEIGHT_0_7037 = 16'd1759;
parameter WEIGHT_0_7038 = 16'd-5641;
parameter WEIGHT_0_7039 = 16'd-10933;
parameter WEIGHT_0_7040 = 16'd-6216;
parameter WEIGHT_0_7041 = 16'd-8776;
parameter WEIGHT_0_7042 = 16'd-6932;
parameter WEIGHT_0_7043 = 16'd1079;
parameter WEIGHT_0_7044 = 16'd-2653;
parameter WEIGHT_0_7045 = 16'd-265;
parameter WEIGHT_0_7046 = 16'd-2193;
parameter WEIGHT_0_7047 = 16'd5700;
parameter WEIGHT_0_7048 = 16'd-13727;
parameter WEIGHT_0_7049 = 16'd-1644;
parameter WEIGHT_0_7050 = 16'd-13210;
parameter WEIGHT_0_7051 = 16'd-12209;
parameter WEIGHT_0_7052 = 16'd-15141;
parameter WEIGHT_0_7053 = 16'd7402;
parameter WEIGHT_0_7054 = 16'd-4270;
parameter WEIGHT_0_7055 = 16'd-5404;
parameter WEIGHT_0_7056 = 16'd-1112;
parameter WEIGHT_0_7057 = 16'd7373;
parameter WEIGHT_0_7058 = 16'd-13219;
parameter WEIGHT_0_7059 = 16'd8181;
parameter WEIGHT_0_7060 = 16'd-12296;
parameter WEIGHT_0_7061 = 16'd-13959;
parameter WEIGHT_0_7062 = 16'd-9681;
parameter WEIGHT_0_7063 = 16'd7256;
parameter WEIGHT_0_7064 = 16'd-9509;
parameter WEIGHT_0_7065 = 16'd-2501;
parameter WEIGHT_0_7066 = 16'd-7372;
parameter WEIGHT_0_7067 = 16'd5560;
parameter WEIGHT_0_7068 = 16'd-11566;
parameter WEIGHT_0_7069 = 16'd8563;
parameter WEIGHT_0_7070 = 16'd-12413;
parameter WEIGHT_0_7071 = 16'd-19023;
parameter WEIGHT_0_7072 = 16'd-16448;
parameter WEIGHT_0_7073 = 16'd11479;
parameter WEIGHT_0_7074 = 16'd-9056;
parameter WEIGHT_0_7075 = 16'd-1435;
parameter WEIGHT_0_7076 = 16'd-3771;
parameter WEIGHT_0_7077 = 16'd8416;
parameter WEIGHT_0_7078 = 16'd-10498;
parameter WEIGHT_0_7079 = 16'd5930;
parameter WEIGHT_0_7080 = 16'd-14705;
parameter WEIGHT_0_7081 = 16'd-9684;
parameter WEIGHT_0_7082 = 16'd-21327;
parameter WEIGHT_0_7083 = 16'd12574;
parameter WEIGHT_0_7084 = 16'd-10020;
parameter WEIGHT_0_7085 = 16'd-1500;
parameter WEIGHT_0_7086 = 16'd-9137;
parameter WEIGHT_0_7087 = 16'd8002;
parameter WEIGHT_0_7088 = 16'd-10506;
parameter WEIGHT_0_7089 = 16'd5444;
parameter WEIGHT_0_7090 = 16'd-19543;
parameter WEIGHT_0_7091 = 16'd-15261;
parameter WEIGHT_0_7092 = 16'd-22418;
parameter WEIGHT_0_7093 = 16'd14403;
parameter WEIGHT_0_7094 = 16'd-8163;
parameter WEIGHT_0_7095 = 16'd328;
parameter WEIGHT_0_7096 = 16'd-10587;
parameter WEIGHT_0_7097 = 16'd9042;
parameter WEIGHT_0_7098 = 16'd-11405;
parameter WEIGHT_0_7099 = 16'd2755;
parameter WEIGHT_0_7100 = 16'd-17975;
parameter WEIGHT_0_7101 = 16'd-19202;
parameter WEIGHT_0_7102 = 16'd-18075;
parameter WEIGHT_0_7103 = 16'd13593;
parameter WEIGHT_0_7104 = 16'd-6101;
parameter WEIGHT_0_7105 = 16'd2069;
parameter WEIGHT_0_7106 = 16'd-8420;
parameter WEIGHT_0_7107 = 16'd8119;
parameter WEIGHT_0_7108 = 16'd-4698;
parameter WEIGHT_0_7109 = 16'd6209;
parameter WEIGHT_0_7110 = 16'd-19336;
parameter WEIGHT_0_7111 = 16'd-22945;
parameter WEIGHT_0_7112 = 16'd-18069;
parameter WEIGHT_0_7113 = 16'd11537;
parameter WEIGHT_0_7114 = 16'd-9267;
parameter WEIGHT_0_7115 = 16'd4969;
parameter WEIGHT_0_7116 = 16'd-7341;
parameter WEIGHT_0_7117 = 16'd5716;
parameter WEIGHT_0_7118 = 16'd-5936;
parameter WEIGHT_0_7119 = 16'd525;
parameter WEIGHT_0_7120 = 16'd-18226;
parameter WEIGHT_0_7121 = 16'd-16507;
parameter WEIGHT_0_7122 = 16'd-13584;
parameter WEIGHT_0_7123 = 16'd12484;
parameter WEIGHT_0_7124 = 16'd-16503;
parameter WEIGHT_0_7125 = 16'd3890;
parameter WEIGHT_0_7126 = 16'd-6759;
parameter WEIGHT_0_7127 = 16'd5297;
parameter WEIGHT_0_7128 = 16'd-6300;
parameter WEIGHT_0_7129 = 16'd2889;
parameter WEIGHT_0_7130 = 16'd-17315;
parameter WEIGHT_0_7131 = 16'd-12683;
parameter WEIGHT_0_7132 = 16'd-12078;
parameter WEIGHT_0_7133 = 16'd11972;
parameter WEIGHT_0_7134 = 16'd-7989;
parameter WEIGHT_0_7135 = 16'd7567;
parameter WEIGHT_0_7136 = 16'd-12787;
parameter WEIGHT_0_7137 = 16'd7092;
parameter WEIGHT_0_7138 = 16'd-3568;
parameter WEIGHT_0_7139 = 16'd2799;
parameter WEIGHT_0_7140 = 16'd-19512;
parameter WEIGHT_0_7141 = 16'd-16424;
parameter WEIGHT_0_7142 = 16'd-4615;
parameter WEIGHT_0_7143 = 16'd5401;
parameter WEIGHT_0_7144 = 16'd-10320;
parameter WEIGHT_0_7145 = 16'd536;
parameter WEIGHT_0_7146 = 16'd-17090;
parameter WEIGHT_0_7147 = 16'd6516;
parameter WEIGHT_0_7148 = 16'd-4321;
parameter WEIGHT_0_7149 = 16'd3740;
parameter WEIGHT_0_7150 = 16'd-22350;
parameter WEIGHT_0_7151 = 16'd-19077;
parameter WEIGHT_0_7152 = 16'd-2550;
parameter WEIGHT_0_7153 = 16'd2926;
parameter WEIGHT_0_7154 = 16'd-9297;
parameter WEIGHT_0_7155 = 16'd4745;
parameter WEIGHT_0_7156 = 16'd-13217;
parameter WEIGHT_0_7157 = 16'd6153;
parameter WEIGHT_0_7158 = 16'd3222;
parameter WEIGHT_0_7159 = 16'd1470;
parameter WEIGHT_0_7160 = 16'd-23173;
parameter WEIGHT_0_7161 = 16'd-22128;
parameter WEIGHT_0_7162 = 16'd-4825;
parameter WEIGHT_0_7163 = 16'd1203;
parameter WEIGHT_0_7164 = 16'd-10388;
parameter WEIGHT_0_7165 = 16'd5911;
parameter WEIGHT_0_7166 = 16'd-16040;
parameter WEIGHT_0_7167 = 16'd6109;
parameter WEIGHT_0_7168 = 16'd-86;
parameter WEIGHT_0_7169 = 16'd5407;
parameter WEIGHT_0_7170 = 16'd-18155;
parameter WEIGHT_0_7171 = 16'd-21607;
parameter WEIGHT_0_7172 = 16'd-8112;
parameter WEIGHT_0_7173 = 16'd400;
parameter WEIGHT_0_7174 = 16'd-12983;
parameter WEIGHT_0_7175 = 16'd5836;
parameter WEIGHT_0_7176 = 16'd-17505;
parameter WEIGHT_0_7177 = 16'd7425;
parameter WEIGHT_0_7178 = 16'd-627;
parameter WEIGHT_0_7179 = 16'd6618;
parameter WEIGHT_0_7180 = 16'd-16594;
parameter WEIGHT_0_7181 = 16'd-19634;
parameter WEIGHT_0_7182 = 16'd-9472;
parameter WEIGHT_0_7183 = 16'd238;
parameter WEIGHT_0_7184 = 16'd-11009;
parameter WEIGHT_0_7185 = 16'd120;
parameter WEIGHT_0_7186 = 16'd-16969;
parameter WEIGHT_0_7187 = 16'd3091;
parameter WEIGHT_0_7188 = 16'd-748;
parameter WEIGHT_0_7189 = 16'd9307;
parameter WEIGHT_0_7190 = 16'd-18858;
parameter WEIGHT_0_7191 = 16'd-11828;
parameter WEIGHT_0_7192 = 16'd-10493;
parameter WEIGHT_0_7193 = 16'd234;
parameter WEIGHT_0_7194 = 16'd-9821;
parameter WEIGHT_0_7195 = 16'd609;
parameter WEIGHT_0_7196 = 16'd-11194;
parameter WEIGHT_0_7197 = 16'd729;
parameter WEIGHT_0_7198 = 16'd387;
parameter WEIGHT_0_7199 = 16'd11184;
parameter WEIGHT_0_7200 = 16'd-11967;
parameter WEIGHT_0_7201 = 16'd-13827;
parameter WEIGHT_0_7202 = 16'd-8279;
parameter WEIGHT_0_7203 = 16'd-1790;
parameter WEIGHT_0_7204 = 16'd-11449;
parameter WEIGHT_0_7205 = 16'd-2451;
parameter WEIGHT_0_7206 = 16'd-11477;
parameter WEIGHT_0_7207 = 16'd-5793;
parameter WEIGHT_0_7208 = 16'd280;
parameter WEIGHT_0_7209 = 16'd14360;
parameter WEIGHT_0_7210 = 16'd-9850;
parameter WEIGHT_0_7211 = 16'd-5948;
parameter WEIGHT_0_7212 = 16'd-7829;
parameter WEIGHT_0_7213 = 16'd-8031;
parameter WEIGHT_0_7214 = 16'd-7202;
parameter WEIGHT_0_7215 = 16'd3554;
parameter WEIGHT_0_7216 = 16'd-5426;
parameter WEIGHT_0_7217 = 16'd69;
parameter WEIGHT_0_7218 = 16'd-12724;
parameter WEIGHT_0_7219 = 16'd12437;
parameter WEIGHT_0_7220 = 16'd-8927;
parameter WEIGHT_0_7221 = 16'd-7661;
parameter WEIGHT_0_7222 = 16'd-10915;
parameter WEIGHT_0_7223 = 16'd-4562;
parameter WEIGHT_0_7224 = 16'd-6114;
parameter WEIGHT_0_7225 = 16'd4235;
parameter WEIGHT_0_7226 = 16'd-3265;
parameter WEIGHT_0_7227 = 16'd-1303;
parameter WEIGHT_0_7228 = 16'd-16774;
parameter WEIGHT_0_7229 = 16'd2362;
parameter WEIGHT_0_7230 = 16'd-7442;
parameter WEIGHT_0_7231 = 16'd-2525;
parameter WEIGHT_0_7232 = 16'd-11163;
parameter WEIGHT_0_7233 = 16'd-8286;
parameter WEIGHT_0_7234 = 16'd-3545;
parameter WEIGHT_0_7235 = 16'd5197;
parameter WEIGHT_0_7236 = 16'd-5203;
parameter WEIGHT_0_7237 = 16'd-6915;
parameter WEIGHT_0_7238 = 16'd-4020;
parameter WEIGHT_0_7239 = 16'd2447;
parameter WEIGHT_0_7240 = 16'd-4551;
parameter WEIGHT_0_7241 = 16'd928;
parameter WEIGHT_0_7242 = 16'd-6319;
parameter WEIGHT_0_7243 = 16'd-672;
parameter WEIGHT_0_7244 = 16'd-5598;
parameter WEIGHT_0_7245 = 16'd3097;
parameter WEIGHT_0_7246 = 16'd-4652;
parameter WEIGHT_0_7247 = 16'd1562;
parameter WEIGHT_0_7248 = 16'd-4785;
parameter WEIGHT_0_7249 = 16'd1914;
parameter WEIGHT_0_7250 = 16'd1396;
parameter WEIGHT_0_7251 = 16'd-464;
parameter WEIGHT_0_7252 = 16'd3370;
parameter WEIGHT_0_7253 = 16'd-3502;
parameter WEIGHT_0_7254 = 16'd-4763;
parameter WEIGHT_0_7255 = 16'd359;
parameter WEIGHT_0_7256 = 16'd686;
parameter WEIGHT_0_7257 = 16'd-534;
parameter WEIGHT_0_7258 = 16'd-6024;
parameter WEIGHT_0_7259 = 16'd-420;
parameter WEIGHT_0_7260 = 16'd1861;
parameter WEIGHT_0_7261 = 16'd-3906;
parameter WEIGHT_0_7262 = 16'd5346;
parameter WEIGHT_0_7263 = 16'd-3346;
parameter WEIGHT_0_7264 = 16'd-3934;
parameter WEIGHT_0_7265 = 16'd-3869;
parameter WEIGHT_0_7266 = 16'd-1091;
parameter WEIGHT_0_7267 = 16'd-3292;
parameter WEIGHT_0_7268 = 16'd-1956;
parameter WEIGHT_0_7269 = 16'd-3016;
parameter WEIGHT_0_7270 = 16'd-142;
parameter WEIGHT_0_7271 = 16'd-110;
parameter WEIGHT_0_7272 = 16'd-685;
parameter WEIGHT_0_7273 = 16'd-591;
parameter WEIGHT_0_7274 = 16'd-1620;
parameter WEIGHT_0_7275 = 16'd-852;
parameter WEIGHT_0_7276 = 16'd1860;
parameter WEIGHT_0_7277 = 16'd2327;
parameter WEIGHT_0_7278 = 16'd920;
parameter WEIGHT_0_7279 = 16'd2203;
parameter WEIGHT_0_7280 = 16'd1308;
parameter WEIGHT_0_7281 = 16'd43;
parameter WEIGHT_0_7282 = 16'd2701;
parameter WEIGHT_0_7283 = 16'd2625;
parameter WEIGHT_0_7284 = 16'd848;
parameter WEIGHT_0_7285 = 16'd2200;
parameter WEIGHT_0_7286 = 16'd1550;
parameter WEIGHT_0_7287 = 16'd446;
parameter WEIGHT_0_7288 = 16'd-395;
parameter WEIGHT_0_7289 = 16'd-1931;
parameter WEIGHT_0_7290 = 16'd2740;
parameter WEIGHT_0_7291 = 16'd-2090;
parameter WEIGHT_0_7292 = 16'd539;
parameter WEIGHT_0_7293 = 16'd680;
parameter WEIGHT_0_7294 = 16'd1179;
parameter WEIGHT_0_7295 = 16'd-1179;
parameter WEIGHT_0_7296 = 16'd1170;
parameter WEIGHT_0_7297 = 16'd2680;
parameter WEIGHT_0_7298 = 16'd676;
parameter WEIGHT_0_7299 = 16'd-564;
parameter WEIGHT_0_7300 = 16'd-419;
parameter WEIGHT_0_7301 = 16'd1319;
parameter WEIGHT_0_7302 = 16'd231;
parameter WEIGHT_0_7303 = 16'd483;
parameter WEIGHT_0_7304 = 16'd-2583;
parameter WEIGHT_0_7305 = 16'd720;
parameter WEIGHT_0_7306 = 16'd-2064;
parameter WEIGHT_0_7307 = 16'd1485;
parameter WEIGHT_0_7308 = 16'd1384;
parameter WEIGHT_0_7309 = 16'd216;
parameter WEIGHT_0_7310 = 16'd-3231;
parameter WEIGHT_0_7311 = 16'd-4120;
parameter WEIGHT_0_7312 = 16'd-2937;
parameter WEIGHT_0_7313 = 16'd-2466;
parameter WEIGHT_0_7314 = 16'd-1874;
parameter WEIGHT_0_7315 = 16'd336;
parameter WEIGHT_0_7316 = 16'd-2993;
parameter WEIGHT_0_7317 = 16'd-1253;
parameter WEIGHT_0_7318 = 16'd261;
parameter WEIGHT_0_7319 = 16'd2275;
parameter WEIGHT_0_7320 = 16'd-2045;
parameter WEIGHT_0_7321 = 16'd-7378;
parameter WEIGHT_0_7322 = 16'd-7277;
parameter WEIGHT_0_7323 = 16'd-4587;
parameter WEIGHT_0_7324 = 16'd-3869;
parameter WEIGHT_0_7325 = 16'd-3990;
parameter WEIGHT_0_7326 = 16'd-1756;
parameter WEIGHT_0_7327 = 16'd-6974;
parameter WEIGHT_0_7328 = 16'd-4530;
parameter WEIGHT_0_7329 = 16'd6389;
parameter WEIGHT_0_7330 = 16'd-6571;
parameter WEIGHT_0_7331 = 16'd-9888;
parameter WEIGHT_0_7332 = 16'd-6178;
parameter WEIGHT_0_7333 = 16'd496;
parameter WEIGHT_0_7334 = 16'd-290;
parameter WEIGHT_0_7335 = 16'd-6791;
parameter WEIGHT_0_7336 = 16'd911;
parameter WEIGHT_0_7337 = 16'd-2839;
parameter WEIGHT_0_7338 = 16'd-5655;
parameter WEIGHT_0_7339 = 16'd7963;
parameter WEIGHT_0_7340 = 16'd-5388;
parameter WEIGHT_0_7341 = 16'd-9693;
parameter WEIGHT_0_7342 = 16'd-6447;
parameter WEIGHT_0_7343 = 16'd-2524;
parameter WEIGHT_0_7344 = 16'd-4011;
parameter WEIGHT_0_7345 = 16'd-11566;
parameter WEIGHT_0_7346 = 16'd67;
parameter WEIGHT_0_7347 = 16'd-3555;
parameter WEIGHT_0_7348 = 16'd-12988;
parameter WEIGHT_0_7349 = 16'd12406;
parameter WEIGHT_0_7350 = 16'd-7538;
parameter WEIGHT_0_7351 = 16'd-7555;
parameter WEIGHT_0_7352 = 16'd-12204;
parameter WEIGHT_0_7353 = 16'd96;
parameter WEIGHT_0_7354 = 16'd-15328;
parameter WEIGHT_0_7355 = 16'd-10984;
parameter WEIGHT_0_7356 = 16'd-2249;
parameter WEIGHT_0_7357 = 16'd70;
parameter WEIGHT_0_7358 = 16'd-9121;
parameter WEIGHT_0_7359 = 16'd7423;
parameter WEIGHT_0_7360 = 16'd-11706;
parameter WEIGHT_0_7361 = 16'd-7061;
parameter WEIGHT_0_7362 = 16'd-12952;
parameter WEIGHT_0_7363 = 16'd-1186;
parameter WEIGHT_0_7364 = 16'd-15979;
parameter WEIGHT_0_7365 = 16'd-8562;
parameter WEIGHT_0_7366 = 16'd-4084;
parameter WEIGHT_0_7367 = 16'd4857;
parameter WEIGHT_0_7368 = 16'd-7003;
parameter WEIGHT_0_7369 = 16'd10160;
parameter WEIGHT_0_7370 = 16'd-17540;
parameter WEIGHT_0_7371 = 16'd-13330;
parameter WEIGHT_0_7372 = 16'd-12230;
parameter WEIGHT_0_7373 = 16'd-1924;
parameter WEIGHT_0_7374 = 16'd-25177;
parameter WEIGHT_0_7375 = 16'd-4485;
parameter WEIGHT_0_7376 = 16'd-6179;
parameter WEIGHT_0_7377 = 16'd6022;
parameter WEIGHT_0_7378 = 16'd-10819;
parameter WEIGHT_0_7379 = 16'd7937;
parameter WEIGHT_0_7380 = 16'd-13069;
parameter WEIGHT_0_7381 = 16'd-7938;
parameter WEIGHT_0_7382 = 16'd-12552;
parameter WEIGHT_0_7383 = 16'd-2750;
parameter WEIGHT_0_7384 = 16'd-18005;
parameter WEIGHT_0_7385 = 16'd-3708;
parameter WEIGHT_0_7386 = 16'd-4276;
parameter WEIGHT_0_7387 = 16'd5522;
parameter WEIGHT_0_7388 = 16'd-10467;
parameter WEIGHT_0_7389 = 16'd9567;
parameter WEIGHT_0_7390 = 16'd-12927;
parameter WEIGHT_0_7391 = 16'd-12761;
parameter WEIGHT_0_7392 = 16'd-12675;
parameter WEIGHT_0_7393 = 16'd-5968;
parameter WEIGHT_0_7394 = 16'd-24488;
parameter WEIGHT_0_7395 = 16'd919;
parameter WEIGHT_0_7396 = 16'd-5282;
parameter WEIGHT_0_7397 = 16'd5491;
parameter WEIGHT_0_7398 = 16'd-9540;
parameter WEIGHT_0_7399 = 16'd5798;
parameter WEIGHT_0_7400 = 16'd-13797;
parameter WEIGHT_0_7401 = 16'd-16674;
parameter WEIGHT_0_7402 = 16'd-16264;
parameter WEIGHT_0_7403 = 16'd-3744;
parameter WEIGHT_0_7404 = 16'd-22501;
parameter WEIGHT_0_7405 = 16'd-886;
parameter WEIGHT_0_7406 = 16'd-5188;
parameter WEIGHT_0_7407 = 16'd2160;
parameter WEIGHT_0_7408 = 16'd-12106;
parameter WEIGHT_0_7409 = 16'd8649;
parameter WEIGHT_0_7410 = 16'd-11643;
parameter WEIGHT_0_7411 = 16'd-18313;
parameter WEIGHT_0_7412 = 16'd-15231;
parameter WEIGHT_0_7413 = 16'd-5219;
parameter WEIGHT_0_7414 = 16'd-29855;
parameter WEIGHT_0_7415 = 16'd-2361;
parameter WEIGHT_0_7416 = 16'd-6317;
parameter WEIGHT_0_7417 = 16'd8912;
parameter WEIGHT_0_7418 = 16'd-12550;
parameter WEIGHT_0_7419 = 16'd9676;
parameter WEIGHT_0_7420 = 16'd-15455;
parameter WEIGHT_0_7421 = 16'd-13188;
parameter WEIGHT_0_7422 = 16'd-16812;
parameter WEIGHT_0_7423 = 16'd-5583;
parameter WEIGHT_0_7424 = 16'd-30561;
parameter WEIGHT_0_7425 = 16'd-3596;
parameter WEIGHT_0_7426 = 16'd-7665;
parameter WEIGHT_0_7427 = 16'd7922;
parameter WEIGHT_0_7428 = 16'd-15013;
parameter WEIGHT_0_7429 = 16'd13789;
parameter WEIGHT_0_7430 = 16'd-16657;
parameter WEIGHT_0_7431 = 16'd-6753;
parameter WEIGHT_0_7432 = 16'd-11761;
parameter WEIGHT_0_7433 = 16'd-6300;
parameter WEIGHT_0_7434 = 16'd-23803;
parameter WEIGHT_0_7435 = 16'd-2125;
parameter WEIGHT_0_7436 = 16'd-5406;
parameter WEIGHT_0_7437 = 16'd11123;
parameter WEIGHT_0_7438 = 16'd-23724;
parameter WEIGHT_0_7439 = 16'd6984;
parameter WEIGHT_0_7440 = 16'd-11520;
parameter WEIGHT_0_7441 = 16'd-10960;
parameter WEIGHT_0_7442 = 16'd-10493;
parameter WEIGHT_0_7443 = 16'd-3625;
parameter WEIGHT_0_7444 = 16'd-27185;
parameter WEIGHT_0_7445 = 16'd645;
parameter WEIGHT_0_7446 = 16'd-7050;
parameter WEIGHT_0_7447 = 16'd10416;
parameter WEIGHT_0_7448 = 16'd-22334;
parameter WEIGHT_0_7449 = 16'd6940;
parameter WEIGHT_0_7450 = 16'd-12187;
parameter WEIGHT_0_7451 = 16'd-12868;
parameter WEIGHT_0_7452 = 16'd-11286;
parameter WEIGHT_0_7453 = 16'd-2727;
parameter WEIGHT_0_7454 = 16'd-22587;
parameter WEIGHT_0_7455 = 16'd-4282;
parameter WEIGHT_0_7456 = 16'd-5157;
parameter WEIGHT_0_7457 = 16'd8223;
parameter WEIGHT_0_7458 = 16'd-13646;
parameter WEIGHT_0_7459 = 16'd5393;
parameter WEIGHT_0_7460 = 16'd-10165;
parameter WEIGHT_0_7461 = 16'd-6373;
parameter WEIGHT_0_7462 = 16'd-15622;
parameter WEIGHT_0_7463 = 16'd-3232;
parameter WEIGHT_0_7464 = 16'd-23000;
parameter WEIGHT_0_7465 = 16'd-4554;
parameter WEIGHT_0_7466 = 16'd-7623;
parameter WEIGHT_0_7467 = 16'd7885;
parameter WEIGHT_0_7468 = 16'd-11775;
parameter WEIGHT_0_7469 = 16'd8024;
parameter WEIGHT_0_7470 = 16'd-7736;
parameter WEIGHT_0_7471 = 16'd-6978;
parameter WEIGHT_0_7472 = 16'd-13175;
parameter WEIGHT_0_7473 = 16'd-725;
parameter WEIGHT_0_7474 = 16'd-17045;
parameter WEIGHT_0_7475 = 16'd-5374;
parameter WEIGHT_0_7476 = 16'd-6433;
parameter WEIGHT_0_7477 = 16'd10372;
parameter WEIGHT_0_7478 = 16'd-18795;
parameter WEIGHT_0_7479 = 16'd7708;
parameter WEIGHT_0_7480 = 16'd-7931;
parameter WEIGHT_0_7481 = 16'd-4898;
parameter WEIGHT_0_7482 = 16'd-8103;
parameter WEIGHT_0_7483 = 16'd1178;
parameter WEIGHT_0_7484 = 16'd-20608;
parameter WEIGHT_0_7485 = 16'd-2181;
parameter WEIGHT_0_7486 = 16'd-5964;
parameter WEIGHT_0_7487 = 16'd-1683;
parameter WEIGHT_0_7488 = 16'd-18528;
parameter WEIGHT_0_7489 = 16'd5344;
parameter WEIGHT_0_7490 = 16'd-7131;
parameter WEIGHT_0_7491 = 16'd-4056;
parameter WEIGHT_0_7492 = 16'd-9062;
parameter WEIGHT_0_7493 = 16'd-3573;
parameter WEIGHT_0_7494 = 16'd-13524;
parameter WEIGHT_0_7495 = 16'd1251;
parameter WEIGHT_0_7496 = 16'd-7539;
parameter WEIGHT_0_7497 = 16'd1321;
parameter WEIGHT_0_7498 = 16'd-14751;
parameter WEIGHT_0_7499 = 16'd5688;
parameter WEIGHT_0_7500 = 16'd-3620;
parameter WEIGHT_0_7501 = 16'd-4313;
parameter WEIGHT_0_7502 = 16'd-9248;
parameter WEIGHT_0_7503 = 16'd-3607;
parameter WEIGHT_0_7504 = 16'd-13027;
parameter WEIGHT_0_7505 = 16'd-1091;
parameter WEIGHT_0_7506 = 16'd-5398;
parameter WEIGHT_0_7507 = 16'd5256;
parameter WEIGHT_0_7508 = 16'd-6846;
parameter WEIGHT_0_7509 = 16'd2057;
parameter WEIGHT_0_7510 = 16'd-4971;
parameter WEIGHT_0_7511 = 16'd-2543;
parameter WEIGHT_0_7512 = 16'd-7711;
parameter WEIGHT_0_7513 = 16'd-3180;
parameter WEIGHT_0_7514 = 16'd-4780;
parameter WEIGHT_0_7515 = 16'd-1247;
parameter WEIGHT_0_7516 = 16'd-4826;
parameter WEIGHT_0_7517 = 16'd-2652;
parameter WEIGHT_0_7518 = 16'd1747;
parameter WEIGHT_0_7519 = 16'd701;
parameter WEIGHT_0_7520 = 16'd1144;
parameter WEIGHT_0_7521 = 16'd2270;
parameter WEIGHT_0_7522 = 16'd174;
parameter WEIGHT_0_7523 = 16'd-902;
parameter WEIGHT_0_7524 = 16'd906;
parameter WEIGHT_0_7525 = 16'd1264;
parameter WEIGHT_0_7526 = 16'd-2193;
parameter WEIGHT_0_7527 = 16'd-144;
parameter WEIGHT_0_7528 = 16'd-3306;
parameter WEIGHT_0_7529 = 16'd1869;
parameter WEIGHT_0_7530 = 16'd-2589;
parameter WEIGHT_0_7531 = 16'd2344;
parameter WEIGHT_0_7532 = 16'd1291;
parameter WEIGHT_0_7533 = 16'd617;
parameter WEIGHT_0_7534 = 16'd-1362;
parameter WEIGHT_0_7535 = 16'd1595;
parameter WEIGHT_0_7536 = 16'd-1695;
parameter WEIGHT_0_7537 = 16'd-620;
parameter WEIGHT_0_7538 = 16'd1344;
parameter WEIGHT_0_7539 = 16'd-1375;
parameter WEIGHT_0_7540 = 16'd1783;
parameter WEIGHT_0_7541 = 16'd1735;
parameter WEIGHT_0_7542 = 16'd2776;
parameter WEIGHT_0_7543 = 16'd2681;
parameter WEIGHT_0_7544 = 16'd-1194;
parameter WEIGHT_0_7545 = 16'd414;
parameter WEIGHT_0_7546 = 16'd-2544;
parameter WEIGHT_0_7547 = 16'd2410;
parameter WEIGHT_0_7548 = 16'd-1525;
parameter WEIGHT_0_7549 = 16'd2415;
parameter WEIGHT_0_7550 = 16'd-1486;
parameter WEIGHT_0_7551 = 16'd1958;
parameter WEIGHT_0_7552 = 16'd-1265;
parameter WEIGHT_0_7553 = 16'd-919;
parameter WEIGHT_0_7554 = 16'd-908;
parameter WEIGHT_0_7555 = 16'd2703;
parameter WEIGHT_0_7556 = 16'd-1779;
parameter WEIGHT_0_7557 = 16'd-275;
parameter WEIGHT_0_7558 = 16'd-1468;
parameter WEIGHT_0_7559 = 16'd-339;
parameter WEIGHT_0_7560 = 16'd-1354;
parameter WEIGHT_0_7561 = 16'd-2010;
parameter WEIGHT_0_7562 = 16'd-1904;
parameter WEIGHT_0_7563 = 16'd-1689;
parameter WEIGHT_0_7564 = 16'd1252;
parameter WEIGHT_0_7565 = 16'd-2294;
parameter WEIGHT_0_7566 = 16'd269;
parameter WEIGHT_0_7567 = 16'd-1288;
parameter WEIGHT_0_7568 = 16'd-880;
parameter WEIGHT_0_7569 = 16'd-1997;
parameter WEIGHT_0_7570 = 16'd-1758;
parameter WEIGHT_0_7571 = 16'd-2610;
parameter WEIGHT_0_7572 = 16'd-1374;
parameter WEIGHT_0_7573 = 16'd-785;
parameter WEIGHT_0_7574 = 16'd1438;
parameter WEIGHT_0_7575 = 16'd-1344;
parameter WEIGHT_0_7576 = 16'd-1324;
parameter WEIGHT_0_7577 = 16'd-160;
parameter WEIGHT_0_7578 = 16'd2739;
parameter WEIGHT_0_7579 = 16'd-1060;
parameter WEIGHT_0_7580 = 16'd-765;
parameter WEIGHT_0_7581 = 16'd1465;
parameter WEIGHT_0_7582 = 16'd-2534;
parameter WEIGHT_0_7583 = 16'd-1244;
parameter WEIGHT_0_7584 = 16'd1416;
parameter WEIGHT_0_7585 = 16'd619;
parameter WEIGHT_0_7586 = 16'd-1740;
parameter WEIGHT_0_7587 = 16'd-414;
parameter WEIGHT_0_7588 = 16'd1878;
parameter WEIGHT_0_7589 = 16'd-2596;
parameter WEIGHT_0_7590 = 16'd439;
parameter WEIGHT_0_7591 = 16'd2157;
parameter WEIGHT_0_7592 = 16'd-2393;
parameter WEIGHT_0_7593 = 16'd522;
parameter WEIGHT_0_7594 = 16'd-282;
parameter WEIGHT_0_7595 = 16'd2536;
parameter WEIGHT_0_7596 = 16'd-780;
parameter WEIGHT_0_7597 = 16'd-1572;
parameter WEIGHT_0_7598 = 16'd565;
parameter WEIGHT_0_7599 = 16'd2086;
parameter WEIGHT_0_7600 = 16'd418;
parameter WEIGHT_0_7601 = 16'd160;
parameter WEIGHT_0_7602 = 16'd584;
parameter WEIGHT_0_7603 = 16'd-3600;
parameter WEIGHT_0_7604 = 16'd-609;
parameter WEIGHT_0_7605 = 16'd-920;
parameter WEIGHT_0_7606 = 16'd827;
parameter WEIGHT_0_7607 = 16'd-127;
parameter WEIGHT_0_7608 = 16'd-641;
parameter WEIGHT_0_7609 = 16'd-3338;
parameter WEIGHT_0_7610 = 16'd468;
parameter WEIGHT_0_7611 = 16'd-1118;
parameter WEIGHT_0_7612 = 16'd607;
parameter WEIGHT_0_7613 = 16'd-25;
parameter WEIGHT_0_7614 = 16'd-4040;
parameter WEIGHT_0_7615 = 16'd-641;
parameter WEIGHT_0_7616 = 16'd-1643;
parameter WEIGHT_0_7617 = 16'd5905;
parameter WEIGHT_0_7618 = 16'd1005;
parameter WEIGHT_0_7619 = 16'd-3475;
parameter WEIGHT_0_7620 = 16'd641;
parameter WEIGHT_0_7621 = 16'd1846;
parameter WEIGHT_0_7622 = 16'd-1053;
parameter WEIGHT_0_7623 = 16'd184;
parameter WEIGHT_0_7624 = 16'd-5740;
parameter WEIGHT_0_7625 = 16'd-3905;
parameter WEIGHT_0_7626 = 16'd-2312;
parameter WEIGHT_0_7627 = 16'd4448;
parameter WEIGHT_0_7628 = 16'd-4234;
parameter WEIGHT_0_7629 = 16'd-2899;
parameter WEIGHT_0_7630 = 16'd-1058;
parameter WEIGHT_0_7631 = 16'd-3433;
parameter WEIGHT_0_7632 = 16'd59;
parameter WEIGHT_0_7633 = 16'd501;
parameter WEIGHT_0_7634 = 16'd-2530;
parameter WEIGHT_0_7635 = 16'd-2521;
parameter WEIGHT_0_7636 = 16'd15;
parameter WEIGHT_0_7637 = 16'd2933;
parameter WEIGHT_0_7638 = 16'd-6672;
parameter WEIGHT_0_7639 = 16'd-2098;
parameter WEIGHT_0_7640 = 16'd-1384;
parameter WEIGHT_0_7641 = 16'd-3048;
parameter WEIGHT_0_7642 = 16'd-1511;
parameter WEIGHT_0_7643 = 16'd943;
parameter WEIGHT_0_7644 = 16'd-6792;
parameter WEIGHT_0_7645 = 16'd-2338;
parameter WEIGHT_0_7646 = 16'd-623;
parameter WEIGHT_0_7647 = 16'd1418;
parameter WEIGHT_0_7648 = 16'd-5975;
parameter WEIGHT_0_7649 = 16'd-1925;
parameter WEIGHT_0_7650 = 16'd-1755;
parameter WEIGHT_0_7651 = 16'd-3260;
parameter WEIGHT_0_7652 = 16'd1373;
parameter WEIGHT_0_7653 = 16'd-6376;
parameter WEIGHT_0_7654 = 16'd-7332;
parameter WEIGHT_0_7655 = 16'd-2004;
parameter WEIGHT_0_7656 = 16'd1417;
parameter WEIGHT_0_7657 = 16'd4159;
parameter WEIGHT_0_7658 = 16'd-6497;
parameter WEIGHT_0_7659 = 16'd-768;
parameter WEIGHT_0_7660 = 16'd-4407;
parameter WEIGHT_0_7661 = 16'd-2121;
parameter WEIGHT_0_7662 = 16'd-5979;
parameter WEIGHT_0_7663 = 16'd-8966;
parameter WEIGHT_0_7664 = 16'd-5499;
parameter WEIGHT_0_7665 = 16'd1387;
parameter WEIGHT_0_7666 = 16'd-1139;
parameter WEIGHT_0_7667 = 16'd5709;
parameter WEIGHT_0_7668 = 16'd-4730;
parameter WEIGHT_0_7669 = 16'd-1629;
parameter WEIGHT_0_7670 = 16'd-5012;
parameter WEIGHT_0_7671 = 16'd-681;
parameter WEIGHT_0_7672 = 16'd-1877;
parameter WEIGHT_0_7673 = 16'd-3225;
parameter WEIGHT_0_7674 = 16'd-10485;
parameter WEIGHT_0_7675 = 16'd-1009;
parameter WEIGHT_0_7676 = 16'd-2740;
parameter WEIGHT_0_7677 = 16'd2232;
parameter WEIGHT_0_7678 = 16'd-7987;
parameter WEIGHT_0_7679 = 16'd-1413;
parameter WEIGHT_0_7680 = 16'd-3843;
parameter WEIGHT_0_7681 = 16'd-975;
parameter WEIGHT_0_7682 = 16'd-1080;
parameter WEIGHT_0_7683 = 16'd-6379;
parameter WEIGHT_0_7684 = 16'd-8094;
parameter WEIGHT_0_7685 = 16'd834;
parameter WEIGHT_0_7686 = 16'd-1146;
parameter WEIGHT_0_7687 = 16'd3976;
parameter WEIGHT_0_7688 = 16'd-8616;
parameter WEIGHT_0_7689 = 16'd-3589;
parameter WEIGHT_0_7690 = 16'd-4092;
parameter WEIGHT_0_7691 = 16'd-4996;
parameter WEIGHT_0_7692 = 16'd-2123;
parameter WEIGHT_0_7693 = 16'd-6833;
parameter WEIGHT_0_7694 = 16'd-11310;
parameter WEIGHT_0_7695 = 16'd-6104;
parameter WEIGHT_0_7696 = 16'd-2081;
parameter WEIGHT_0_7697 = 16'd15895;
parameter WEIGHT_0_7698 = 16'd-8260;
parameter WEIGHT_0_7699 = 16'd-9898;
parameter WEIGHT_0_7700 = 16'd-9047;
parameter WEIGHT_0_7701 = 16'd-5947;
parameter WEIGHT_0_7702 = 16'd-1476;
parameter WEIGHT_0_7703 = 16'd-8740;
parameter WEIGHT_0_7704 = 16'd-14965;
parameter WEIGHT_0_7705 = 16'd-9412;
parameter WEIGHT_0_7706 = 16'd-5583;
parameter WEIGHT_0_7707 = 16'd8292;
parameter WEIGHT_0_7708 = 16'd-10094;
parameter WEIGHT_0_7709 = 16'd-3422;
parameter WEIGHT_0_7710 = 16'd-8171;
parameter WEIGHT_0_7711 = 16'd1040;
parameter WEIGHT_0_7712 = 16'd-997;
parameter WEIGHT_0_7713 = 16'd-6448;
parameter WEIGHT_0_7714 = 16'd-9132;
parameter WEIGHT_0_7715 = 16'd-10139;
parameter WEIGHT_0_7716 = 16'd-2643;
parameter WEIGHT_0_7717 = 16'd5011;
parameter WEIGHT_0_7718 = 16'd-4420;
parameter WEIGHT_0_7719 = 16'd-3506;
parameter WEIGHT_0_7720 = 16'd-6759;
parameter WEIGHT_0_7721 = 16'd-1040;
parameter WEIGHT_0_7722 = 16'd672;
parameter WEIGHT_0_7723 = 16'd-9365;
parameter WEIGHT_0_7724 = 16'd-8709;
parameter WEIGHT_0_7725 = 16'd-5893;
parameter WEIGHT_0_7726 = 16'd-1959;
parameter WEIGHT_0_7727 = 16'd8564;
parameter WEIGHT_0_7728 = 16'd-3881;
parameter WEIGHT_0_7729 = 16'd-7100;
parameter WEIGHT_0_7730 = 16'd-4741;
parameter WEIGHT_0_7731 = 16'd-3864;
parameter WEIGHT_0_7732 = 16'd-67;
parameter WEIGHT_0_7733 = 16'd-7968;
parameter WEIGHT_0_7734 = 16'd-9257;
parameter WEIGHT_0_7735 = 16'd-6277;
parameter WEIGHT_0_7736 = 16'd-1682;
parameter WEIGHT_0_7737 = 16'd12251;
parameter WEIGHT_0_7738 = 16'd-5705;
parameter WEIGHT_0_7739 = 16'd-14940;
parameter WEIGHT_0_7740 = 16'd-5741;
parameter WEIGHT_0_7741 = 16'd-5773;
parameter WEIGHT_0_7742 = 16'd-9153;
parameter WEIGHT_0_7743 = 16'd-9757;
parameter WEIGHT_0_7744 = 16'd-8711;
parameter WEIGHT_0_7745 = 16'd-8475;
parameter WEIGHT_0_7746 = 16'd-7210;
parameter WEIGHT_0_7747 = 16'd11281;
parameter WEIGHT_0_7748 = 16'd-11840;
parameter WEIGHT_0_7749 = 16'd-4313;
parameter WEIGHT_0_7750 = 16'd-3584;
parameter WEIGHT_0_7751 = 16'd-3122;
parameter WEIGHT_0_7752 = 16'd-8193;
parameter WEIGHT_0_7753 = 16'd-6294;
parameter WEIGHT_0_7754 = 16'd-4526;
parameter WEIGHT_0_7755 = 16'd-5521;
parameter WEIGHT_0_7756 = 16'd-4503;
parameter WEIGHT_0_7757 = 16'd9167;
parameter WEIGHT_0_7758 = 16'd-6918;
parameter WEIGHT_0_7759 = 16'd-4511;
parameter WEIGHT_0_7760 = 16'd-2055;
parameter WEIGHT_0_7761 = 16'd-1001;
parameter WEIGHT_0_7762 = 16'd-4431;
parameter WEIGHT_0_7763 = 16'd-8830;
parameter WEIGHT_0_7764 = 16'd-2003;
parameter WEIGHT_0_7765 = 16'd-7644;
parameter WEIGHT_0_7766 = 16'd-1432;
parameter WEIGHT_0_7767 = 16'd3392;
parameter WEIGHT_0_7768 = 16'd-5545;
parameter WEIGHT_0_7769 = 16'd2024;
parameter WEIGHT_0_7770 = 16'd-8030;
parameter WEIGHT_0_7771 = 16'd430;
parameter WEIGHT_0_7772 = 16'd-4803;
parameter WEIGHT_0_7773 = 16'd-9451;
parameter WEIGHT_0_7774 = 16'd-5530;
parameter WEIGHT_0_7775 = 16'd-6685;
parameter WEIGHT_0_7776 = 16'd-5042;
parameter WEIGHT_0_7777 = 16'd4381;
parameter WEIGHT_0_7778 = 16'd-10093;
parameter WEIGHT_0_7779 = 16'd8;
parameter WEIGHT_0_7780 = 16'd-6669;
parameter WEIGHT_0_7781 = 16'd-4935;
parameter WEIGHT_0_7782 = 16'd-6806;
parameter WEIGHT_0_7783 = 16'd-4083;
parameter WEIGHT_0_7784 = 16'd-3171;
parameter WEIGHT_0_7785 = 16'd-3076;
parameter WEIGHT_0_7786 = 16'd-2166;
parameter WEIGHT_0_7787 = 16'd4425;
parameter WEIGHT_0_7788 = 16'd-2719;
parameter WEIGHT_0_7789 = 16'd-2399;
parameter WEIGHT_0_7790 = 16'd-2072;
parameter WEIGHT_0_7791 = 16'd591;
parameter WEIGHT_0_7792 = 16'd-3596;
parameter WEIGHT_0_7793 = 16'd-3663;
parameter WEIGHT_0_7794 = 16'd-7123;
parameter WEIGHT_0_7795 = 16'd-2251;
parameter WEIGHT_0_7796 = 16'd-1034;
parameter WEIGHT_0_7797 = 16'd3943;
parameter WEIGHT_0_7798 = 16'd-4536;
parameter WEIGHT_0_7799 = 16'd-6439;
parameter WEIGHT_0_7800 = 16'd-22;
parameter WEIGHT_0_7801 = 16'd-403;
parameter WEIGHT_0_7802 = 16'd2035;
parameter WEIGHT_0_7803 = 16'd-60;
parameter WEIGHT_0_7804 = 16'd-800;
parameter WEIGHT_0_7805 = 16'd1612;
parameter WEIGHT_0_7806 = 16'd2427;
parameter WEIGHT_0_7807 = 16'd2772;
parameter WEIGHT_0_7808 = 16'd2238;
parameter WEIGHT_0_7809 = 16'd17;
parameter WEIGHT_0_7810 = 16'd-2805;
parameter WEIGHT_0_7811 = 16'd-594;
parameter WEIGHT_0_7812 = 16'd-1551;
parameter WEIGHT_0_7813 = 16'd2368;
parameter WEIGHT_0_7814 = 16'd671;
parameter WEIGHT_0_7815 = 16'd1941;
parameter WEIGHT_0_7816 = 16'd-2133;
parameter WEIGHT_0_7817 = 16'd-558;
parameter WEIGHT_0_7818 = 16'd-169;
parameter WEIGHT_0_7819 = 16'd-2585;
parameter WEIGHT_0_7820 = 16'd382;
parameter WEIGHT_0_7821 = 16'd2741;
parameter WEIGHT_0_7822 = 16'd-2706;
parameter WEIGHT_0_7823 = 16'd84;
parameter WEIGHT_0_7824 = 16'd2598;
parameter WEIGHT_0_7825 = 16'd-205;
parameter WEIGHT_0_7826 = 16'd-1950;
parameter WEIGHT_0_7827 = 16'd-531;
parameter WEIGHT_0_7828 = 16'd-567;
parameter WEIGHT_0_7829 = 16'd-376;
parameter WEIGHT_0_7830 = 16'd2362;
parameter WEIGHT_0_7831 = 16'd2501;
parameter WEIGHT_0_7832 = 16'd-729;
parameter WEIGHT_0_7833 = 16'd604;
parameter WEIGHT_0_7834 = 16'd639;
parameter WEIGHT_0_7835 = 16'd1439;
parameter WEIGHT_0_7836 = 16'd-1496;
parameter WEIGHT_0_7837 = 16'd-285;
parameter WEIGHT_0_7838 = 16'd163;
parameter WEIGHT_0_7839 = 16'd-1452;
parameter BIAS_0 = 16'd[ -9078  12758   1249  -6335   2787  19507  -2379  12007 -24979  -4115];

endmodule